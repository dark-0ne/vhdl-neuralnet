----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    20:49:00 02/02/2019 
-- Design Name: 
-- Module Name:    sigmoid - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity sigmoid is
    Port ( Y : in  STD_LOGIC_VECTOR (15 downto 0);
           O : out  STD_LOGIC_VECTOR (15 downto 0));
end sigmoid;

architecture Behavioral of sigmoid is
    type rom is array (0 to 65535) of STD_LOGIC_VECTOR (15 downto 0);
    signal sigmoid_val : rom := (x"07ff", x"07ff", x"07ff", x"0800", x"0800", x"0800", x"0800", x"0801", x"0801", x"0801", x"0801", x"0802", x"0802", x"0802", x"0802", x"0803", x"0803", x"0803", x"0803", x"0804", x"0804", x"0804", x"0804", x"0805", x"0805", x"0805", x"0805", x"0806", x"0806", x"0806", x"0806", x"0807", x"0807", x"0807", x"0807", x"0808", x"0808", x"0808", x"0808", x"0809", x"0809", x"0809", x"0809", x"080a", x"080a", x"080a", x"080a", x"080b", x"080b", x"080b", x"080b", x"080c", x"080c", x"080c", x"080c", x"080d", x"080d", x"080d", x"080d", x"080e", x"080e", x"080e", x"080e", x"080f", x"080f", x"080f", x"080f", x"0810", x"0810", x"0810", x"0810", x"0811", x"0811", x"0811", x"0811", x"0812", x"0812", x"0812", x"0812", x"0813", x"0813", x"0813", x"0813", x"0814", x"0814", x"0814", x"0814", x"0815", x"0815", x"0815", x"0815", x"0816", x"0816", x"0816", x"0816", x"0817", x"0817", x"0817", x"0817", x"0818", x"0818", x"0818", x"0818", x"0819", x"0819", x"0819", x"0819", x"081a", x"081a", x"081a", x"081a", x"081b", x"081b", x"081b", x"081b", x"081c", x"081c", x"081c", x"081c", x"081d", x"081d", x"081d", x"081d", x"081e", x"081e", x"081e", x"081e", x"081f", x"081f", x"081f", x"081f", x"0820", x"0820", x"0820", x"0820", x"0821", x"0821", x"0821", x"0821", x"0822", x"0822", x"0822", x"0822", x"0823", x"0823", x"0823", x"0823", x"0824", x"0824", x"0824", x"0824", x"0825", x"0825", x"0825", x"0825", x"0826", x"0826", x"0826", x"0826", x"0827", x"0827", x"0827", x"0827", x"0828", x"0828", x"0828", x"0828", x"0829", x"0829", x"0829", x"0829", x"082a", x"082a", x"082a", x"082a", x"082b", x"082b", x"082b", x"082b", x"082c", x"082c", x"082c", x"082c", x"082d", x"082d", x"082d", x"082d", x"082e", x"082e", x"082e", x"082e", x"082f", x"082f", x"082f", x"082f", x"0830", x"0830", x"0830", x"0830", x"0831", x"0831", x"0831", x"0831", x"0832", x"0832", x"0832", x"0832", x"0833", x"0833", x"0833", x"0833", x"0834", x"0834", x"0834", x"0834", x"0835", x"0835", x"0835", x"0835", x"0836", x"0836", x"0836", x"0836", x"0837", x"0837", x"0837", x"0837", x"0838", x"0838", x"0838", x"0838", x"0839", x"0839", x"0839", x"0839", x"083a", x"083a", x"083a", x"083a", x"083b", x"083b", x"083b", x"083b", x"083c", x"083c", x"083c", x"083c", x"083d", x"083d", x"083d", x"083d", x"083e", x"083e", x"083e", x"083e", x"083f", x"083f", x"083f", x"083f", x"0840", x"0840", x"0840", x"0840", x"0841", x"0841", x"0841", x"0841", x"0842", x"0842", x"0842", x"0842", x"0843", x"0843", x"0843", x"0843", x"0844", x"0844", x"0844", x"0844", x"0845", x"0845", x"0845", x"0845", x"0846", x"0846", x"0846", x"0846", x"0847", x"0847", x"0847", x"0847", x"0848", x"0848", x"0848", x"0848", x"0849", x"0849", x"0849", x"0849", x"084a", x"084a", x"084a", x"084a", x"084b", x"084b", x"084b", x"084b", x"084c", x"084c", x"084c", x"084c", x"084d", x"084d", x"084d", x"084d", x"084e", x"084e", x"084e", x"084e", x"084f", x"084f", x"084f", x"084f", x"0850", x"0850", x"0850", x"0850", x"0851", x"0851", x"0851", x"0851", x"0852", x"0852", x"0852", x"0852", x"0853", x"0853", x"0853", x"0853", x"0854", x"0854", x"0854", x"0854", x"0855", x"0855", x"0855", x"0855", x"0856", x"0856", x"0856", x"0856", x"0857", x"0857", x"0857", x"0857", x"0858", x"0858", x"0858", x"0858", x"0859", x"0859", x"0859", x"0859", x"085a", x"085a", x"085a", x"085a", x"085b", x"085b", x"085b", x"085b", x"085c", x"085c", x"085c", x"085c", x"085d", x"085d", x"085d", x"085d", x"085e", x"085e", x"085e", x"085e", x"085f", x"085f", x"085f", x"085f", x"0860", x"0860", x"0860", x"0860", x"0861", x"0861", x"0861", x"0861", x"0862", x"0862", x"0862", x"0862", x"0863", x"0863", x"0863", x"0863", x"0864", x"0864", x"0864", x"0864", x"0865", x"0865", x"0865", x"0865", x"0866", x"0866", x"0866", x"0866", x"0867", x"0867", x"0867", x"0867", x"0868", x"0868", x"0868", x"0868", x"0869", x"0869", x"0869", x"0869", x"086a", x"086a", x"086a", x"086a", x"086b", x"086b", x"086b", x"086b", x"086c", x"086c", x"086c", x"086c", x"086d", x"086d", x"086d", x"086d", x"086e", x"086e", x"086e", x"086e", x"086f", x"086f", x"086f", x"086f", x"0870", x"0870", x"0870", x"0870", x"0871", x"0871", x"0871", x"0871", x"0872", x"0872", x"0872", x"0872", x"0873", x"0873", x"0873", x"0873", x"0874", x"0874", x"0874", x"0874", x"0875", x"0875", x"0875", x"0875", x"0876", x"0876", x"0876", x"0876", x"0877", x"0877", x"0877", x"0877", x"0878", x"0878", x"0878", x"0878", x"0879", x"0879", x"0879", x"0879", x"087a", x"087a", x"087a", x"087a", x"087b", x"087b", x"087b", x"087b", x"087c", x"087c", x"087c", x"087c", x"087d", x"087d", x"087d", x"087d", x"087e", x"087e", x"087e", x"087e", x"087f", x"087f", x"087f", x"087f", x"0880", x"0880", x"0880", x"0880", x"0881", x"0881", x"0881", x"0881", x"0882", x"0882", x"0882", x"0882", x"0883", x"0883", x"0883", x"0883", x"0884", x"0884", x"0884", x"0884", x"0885", x"0885", x"0885", x"0885", x"0886", x"0886", x"0886", x"0886", x"0887", x"0887", x"0887", x"0887", x"0888", x"0888", x"0888", x"0888", x"0889", x"0889", x"0889", x"0889", x"088a", x"088a", x"088a", x"088a", x"088a", x"088b", x"088b", x"088b", x"088b", x"088c", x"088c", x"088c", x"088c", x"088d", x"088d", x"088d", x"088d", x"088e", x"088e", x"088e", x"088e", x"088f", x"088f", x"088f", x"088f", x"0890", x"0890", x"0890", x"0890", x"0891", x"0891", x"0891", x"0891", x"0892", x"0892", x"0892", x"0892", x"0893", x"0893", x"0893", x"0893", x"0894", x"0894", x"0894", x"0894", x"0895", x"0895", x"0895", x"0895", x"0896", x"0896", x"0896", x"0896", x"0897", x"0897", x"0897", x"0897", x"0898", x"0898", x"0898", x"0898", x"0899", x"0899", x"0899", x"0899", x"089a", x"089a", x"089a", x"089a", x"089b", x"089b", x"089b", x"089b", x"089c", x"089c", x"089c", x"089c", x"089d", x"089d", x"089d", x"089d", x"089e", x"089e", x"089e", x"089e", x"089f", x"089f", x"089f", x"089f", x"08a0", x"08a0", x"08a0", x"08a0", x"08a1", x"08a1", x"08a1", x"08a1", x"08a2", x"08a2", x"08a2", x"08a2", x"08a3", x"08a3", x"08a3", x"08a3", x"08a4", x"08a4", x"08a4", x"08a4", x"08a5", x"08a5", x"08a5", x"08a5", x"08a6", x"08a6", x"08a6", x"08a6", x"08a7", x"08a7", x"08a7", x"08a7", x"08a8", x"08a8", x"08a8", x"08a8", x"08a9", x"08a9", x"08a9", x"08a9", x"08aa", x"08aa", x"08aa", x"08aa", x"08ab", x"08ab", x"08ab", x"08ab", x"08ac", x"08ac", x"08ac", x"08ac", x"08ad", x"08ad", x"08ad", x"08ad", x"08ae", x"08ae", x"08ae", x"08ae", x"08af", x"08af", x"08af", x"08af", x"08b0", x"08b0", x"08b0", x"08b0", x"08b1", x"08b1", x"08b1", x"08b1", x"08b2", x"08b2", x"08b2", x"08b2", x"08b2", x"08b3", x"08b3", x"08b3", x"08b3", x"08b4", x"08b4", x"08b4", x"08b4", x"08b5", x"08b5", x"08b5", x"08b5", x"08b6", x"08b6", x"08b6", x"08b6", x"08b7", x"08b7", x"08b7", x"08b7", x"08b8", x"08b8", x"08b8", x"08b8", x"08b9", x"08b9", x"08b9", x"08b9", x"08ba", x"08ba", x"08ba", x"08ba", x"08bb", x"08bb", x"08bb", x"08bb", x"08bc", x"08bc", x"08bc", x"08bc", x"08bd", x"08bd", x"08bd", x"08bd", x"08be", x"08be", x"08be", x"08be", x"08bf", x"08bf", x"08bf", x"08bf", x"08c0", x"08c0", x"08c0", x"08c0", x"08c1", x"08c1", x"08c1", x"08c1", x"08c2", x"08c2", x"08c2", x"08c2", x"08c3", x"08c3", x"08c3", x"08c3", x"08c4", x"08c4", x"08c4", x"08c4", x"08c5", x"08c5", x"08c5", x"08c5", x"08c6", x"08c6", x"08c6", x"08c6", x"08c7", x"08c7", x"08c7", x"08c7", x"08c8", x"08c8", x"08c8", x"08c8", x"08c9", x"08c9", x"08c9", x"08c9", x"08ca", x"08ca", x"08ca", x"08ca", x"08cb", x"08cb", x"08cb", x"08cb", x"08cc", x"08cc", x"08cc", x"08cc", x"08cd", x"08cd", x"08cd", x"08cd", x"08cd", x"08ce", x"08ce", x"08ce", x"08ce", x"08cf", x"08cf", x"08cf", x"08cf", x"08d0", x"08d0", x"08d0", x"08d0", x"08d1", x"08d1", x"08d1", x"08d1", x"08d2", x"08d2", x"08d2", x"08d2", x"08d3", x"08d3", x"08d3", x"08d3", x"08d4", x"08d4", x"08d4", x"08d4", x"08d5", x"08d5", x"08d5", x"08d5", x"08d6", x"08d6", x"08d6", x"08d6", x"08d7", x"08d7", x"08d7", x"08d7", x"08d8", x"08d8", x"08d8", x"08d8", x"08d9", x"08d9", x"08d9", x"08d9", x"08da", x"08da", x"08da", x"08da", x"08db", x"08db", x"08db", x"08db", x"08dc", x"08dc", x"08dc", x"08dc", x"08dd", x"08dd", x"08dd", x"08dd", x"08de", x"08de", x"08de", x"08de", x"08df", x"08df", x"08df", x"08df", x"08e0", x"08e0", x"08e0", x"08e0", x"08e1", x"08e1", x"08e1", x"08e1", x"08e2", x"08e2", x"08e2", x"08e2", x"08e3", x"08e3", x"08e3", x"08e3", x"08e3", x"08e4", x"08e4", x"08e4", x"08e4", x"08e5", x"08e5", x"08e5", x"08e5", x"08e6", x"08e6", x"08e6", x"08e6", x"08e7", x"08e7", x"08e7", x"08e7", x"08e8", x"08e8", x"08e8", x"08e8", x"08e9", x"08e9", x"08e9", x"08e9", x"08ea", x"08ea", x"08ea", x"08ea", x"08eb", x"08eb", x"08eb", x"08eb", x"08ec", x"08ec", x"08ec", x"08ec", x"08ed", x"08ed", x"08ed", x"08ed", x"08ee", x"08ee", x"08ee", x"08ee", x"08ef", x"08ef", x"08ef", x"08ef", x"08f0", x"08f0", x"08f0", x"08f0", x"08f1", x"08f1", x"08f1", x"08f1", x"08f2", x"08f2", x"08f2", x"08f2", x"08f3", x"08f3", x"08f3", x"08f3", x"08f4", x"08f4", x"08f4", x"08f4", x"08f5", x"08f5", x"08f5", x"08f5", x"08f5", x"08f6", x"08f6", x"08f6", x"08f6", x"08f7", x"08f7", x"08f7", x"08f7", x"08f8", x"08f8", x"08f8", x"08f8", x"08f9", x"08f9", x"08f9", x"08f9", x"08fa", x"08fa", x"08fa", x"08fa", x"08fb", x"08fb", x"08fb", x"08fb", x"08fc", x"08fc", x"08fc", x"08fc", x"08fd", x"08fd", x"08fd", x"08fd", x"08fe", x"08fe", x"08fe", x"08fe", x"08ff", x"08ff", x"08ff", x"08ff", x"0900", x"0900", x"0900", x"0900", x"0901", x"0901", x"0901", x"0901", x"0902", x"0902", x"0902", x"0902", x"0903", x"0903", x"0903", x"0903", x"0904", x"0904", x"0904", x"0904", x"0904", x"0905", x"0905", x"0905", x"0905", x"0906", x"0906", x"0906", x"0906", x"0907", x"0907", x"0907", x"0907", x"0908", x"0908", x"0908", x"0908", x"0909", x"0909", x"0909", x"0909", x"090a", x"090a", x"090a", x"090a", x"090b", x"090b", x"090b", x"090b", x"090c", x"090c", x"090c", x"090c", x"090d", x"090d", x"090d", x"090d", x"090e", x"090e", x"090e", x"090e", x"090f", x"090f", x"090f", x"090f", x"0910", x"0910", x"0910", x"0910", x"0911", x"0911", x"0911", x"0911", x"0912", x"0912", x"0912", x"0912", x"0913", x"0913", x"0913", x"0913", x"0913", x"0914", x"0914", x"0914", x"0914", x"0915", x"0915", x"0915", x"0915", x"0916", x"0916", x"0916", x"0916", x"0917", x"0917", x"0917", x"0917", x"0918", x"0918", x"0918", x"0918", x"0919", x"0919", x"0919", x"0919", x"091a", x"091a", x"091a", x"091a", x"091b", x"091b", x"091b", x"091b", x"091c", x"091c", x"091c", x"091c", x"091d", x"091d", x"091d", x"091d", x"091e", x"091e", x"091e", x"091e", x"091f", x"091f", x"091f", x"091f", x"091f", x"0920", x"0920", x"0920", x"0920", x"0921", x"0921", x"0921", x"0921", x"0922", x"0922", x"0922", x"0922", x"0923", x"0923", x"0923", x"0923", x"0924", x"0924", x"0924", x"0924", x"0925", x"0925", x"0925", x"0925", x"0926", x"0926", x"0926", x"0926", x"0927", x"0927", x"0927", x"0927", x"0928", x"0928", x"0928", x"0928", x"0929", x"0929", x"0929", x"0929", x"092a", x"092a", x"092a", x"092a", x"092b", x"092b", x"092b", x"092b", x"092b", x"092c", x"092c", x"092c", x"092c", x"092d", x"092d", x"092d", x"092d", x"092e", x"092e", x"092e", x"092e", x"092f", x"092f", x"092f", x"092f", x"0930", x"0930", x"0930", x"0930", x"0931", x"0931", x"0931", x"0931", x"0932", x"0932", x"0932", x"0932", x"0933", x"0933", x"0933", x"0933", x"0934", x"0934", x"0934", x"0934", x"0935", x"0935", x"0935", x"0935", x"0936", x"0936", x"0936", x"0936", x"0936", x"0937", x"0937", x"0937", x"0937", x"0938", x"0938", x"0938", x"0938", x"0939", x"0939", x"0939", x"0939", x"093a", x"093a", x"093a", x"093a", x"093b", x"093b", x"093b", x"093b", x"093c", x"093c", x"093c", x"093c", x"093d", x"093d", x"093d", x"093d", x"093e", x"093e", x"093e", x"093e", x"093f", x"093f", x"093f", x"093f", x"0940", x"0940", x"0940", x"0940", x"0940", x"0941", x"0941", x"0941", x"0941", x"0942", x"0942", x"0942", x"0942", x"0943", x"0943", x"0943", x"0943", x"0944", x"0944", x"0944", x"0944", x"0945", x"0945", x"0945", x"0945", x"0946", x"0946", x"0946", x"0946", x"0947", x"0947", x"0947", x"0947", x"0948", x"0948", x"0948", x"0948", x"0949", x"0949", x"0949", x"0949", x"094a", x"094a", x"094a", x"094a", x"094a", x"094b", x"094b", x"094b", x"094b", x"094c", x"094c", x"094c", x"094c", x"094d", x"094d", x"094d", x"094d", x"094e", x"094e", x"094e", x"094e", x"094f", x"094f", x"094f", x"094f", x"0950", x"0950", x"0950", x"0950", x"0951", x"0951", x"0951", x"0951", x"0952", x"0952", x"0952", x"0952", x"0953", x"0953", x"0953", x"0953", x"0953", x"0954", x"0954", x"0954", x"0954", x"0955", x"0955", x"0955", x"0955", x"0956", x"0956", x"0956", x"0956", x"0957", x"0957", x"0957", x"0957", x"0958", x"0958", x"0958", x"0958", x"0959", x"0959", x"0959", x"0959", x"095a", x"095a", x"095a", x"095a", x"095b", x"095b", x"095b", x"095b", x"095b", x"095c", x"095c", x"095c", x"095c", x"095d", x"095d", x"095d", x"095d", x"095e", x"095e", x"095e", x"095e", x"095f", x"095f", x"095f", x"095f", x"0960", x"0960", x"0960", x"0960", x"0961", x"0961", x"0961", x"0961", x"0962", x"0962", x"0962", x"0962", x"0963", x"0963", x"0963", x"0963", x"0963", x"0964", x"0964", x"0964", x"0964", x"0965", x"0965", x"0965", x"0965", x"0966", x"0966", x"0966", x"0966", x"0967", x"0967", x"0967", x"0967", x"0968", x"0968", x"0968", x"0968", x"0969", x"0969", x"0969", x"0969", x"096a", x"096a", x"096a", x"096a", x"096b", x"096b", x"096b", x"096b", x"096b", x"096c", x"096c", x"096c", x"096c", x"096d", x"096d", x"096d", x"096d", x"096e", x"096e", x"096e", x"096e", x"096f", x"096f", x"096f", x"096f", x"0970", x"0970", x"0970", x"0970", x"0971", x"0971", x"0971", x"0971", x"0972", x"0972", x"0972", x"0972", x"0972", x"0973", x"0973", x"0973", x"0973", x"0974", x"0974", x"0974", x"0974", x"0975", x"0975", x"0975", x"0975", x"0976", x"0976", x"0976", x"0976", x"0977", x"0977", x"0977", x"0977", x"0978", x"0978", x"0978", x"0978", x"0979", x"0979", x"0979", x"0979", x"097a", x"097a", x"097a", x"097a", x"097a", x"097b", x"097b", x"097b", x"097b", x"097c", x"097c", x"097c", x"097c", x"097d", x"097d", x"097d", x"097d", x"097e", x"097e", x"097e", x"097e", x"097f", x"097f", x"097f", x"097f", x"0980", x"0980", x"0980", x"0980", x"0981", x"0981", x"0981", x"0981", x"0981", x"0982", x"0982", x"0982", x"0982", x"0983", x"0983", x"0983", x"0983", x"0984", x"0984", x"0984", x"0984", x"0985", x"0985", x"0985", x"0985", x"0986", x"0986", x"0986", x"0986", x"0987", x"0987", x"0987", x"0987", x"0987", x"0988", x"0988", x"0988", x"0988", x"0989", x"0989", x"0989", x"0989", x"098a", x"098a", x"098a", x"098a", x"098b", x"098b", x"098b", x"098b", x"098c", x"098c", x"098c", x"098c", x"098d", x"098d", x"098d", x"098d", x"098e", x"098e", x"098e", x"098e", x"098e", x"098f", x"098f", x"098f", x"098f", x"0990", x"0990", x"0990", x"0990", x"0991", x"0991", x"0991", x"0991", x"0992", x"0992", x"0992", x"0992", x"0993", x"0993", x"0993", x"0993", x"0994", x"0994", x"0994", x"0994", x"0994", x"0995", x"0995", x"0995", x"0995", x"0996", x"0996", x"0996", x"0996", x"0997", x"0997", x"0997", x"0997", x"0998", x"0998", x"0998", x"0998", x"0999", x"0999", x"0999", x"0999", x"099a", x"099a", x"099a", x"099a", x"099a", x"099b", x"099b", x"099b", x"099b", x"099c", x"099c", x"099c", x"099c", x"099d", x"099d", x"099d", x"099d", x"099e", x"099e", x"099e", x"099e", x"099f", x"099f", x"099f", x"099f", x"09a0", x"09a0", x"09a0", x"09a0", x"09a0", x"09a1", x"09a1", x"09a1", x"09a1", x"09a2", x"09a2", x"09a2", x"09a2", x"09a3", x"09a3", x"09a3", x"09a3", x"09a4", x"09a4", x"09a4", x"09a4", x"09a5", x"09a5", x"09a5", x"09a5", x"09a5", x"09a6", x"09a6", x"09a6", x"09a6", x"09a7", x"09a7", x"09a7", x"09a7", x"09a8", x"09a8", x"09a8", x"09a8", x"09a9", x"09a9", x"09a9", x"09a9", x"09aa", x"09aa", x"09aa", x"09aa", x"09ab", x"09ab", x"09ab", x"09ab", x"09ab", x"09ac", x"09ac", x"09ac", x"09ac", x"09ad", x"09ad", x"09ad", x"09ad", x"09ae", x"09ae", x"09ae", x"09ae", x"09af", x"09af", x"09af", x"09af", x"09b0", x"09b0", x"09b0", x"09b0", x"09b0", x"09b1", x"09b1", x"09b1", x"09b1", x"09b2", x"09b2", x"09b2", x"09b2", x"09b3", x"09b3", x"09b3", x"09b3", x"09b4", x"09b4", x"09b4", x"09b4", x"09b5", x"09b5", x"09b5", x"09b5", x"09b5", x"09b6", x"09b6", x"09b6", x"09b6", x"09b7", x"09b7", x"09b7", x"09b7", x"09b8", x"09b8", x"09b8", x"09b8", x"09b9", x"09b9", x"09b9", x"09b9", x"09ba", x"09ba", x"09ba", x"09ba", x"09bb", x"09bb", x"09bb", x"09bb", x"09bb", x"09bc", x"09bc", x"09bc", x"09bc", x"09bd", x"09bd", x"09bd", x"09bd", x"09be", x"09be", x"09be", x"09be", x"09bf", x"09bf", x"09bf", x"09bf", x"09c0", x"09c0", x"09c0", x"09c0", x"09c0", x"09c1", x"09c1", x"09c1", x"09c1", x"09c2", x"09c2", x"09c2", x"09c2", x"09c3", x"09c3", x"09c3", x"09c3", x"09c4", x"09c4", x"09c4", x"09c4", x"09c4", x"09c5", x"09c5", x"09c5", x"09c5", x"09c6", x"09c6", x"09c6", x"09c6", x"09c7", x"09c7", x"09c7", x"09c7", x"09c8", x"09c8", x"09c8", x"09c8", x"09c9", x"09c9", x"09c9", x"09c9", x"09c9", x"09ca", x"09ca", x"09ca", x"09ca", x"09cb", x"09cb", x"09cb", x"09cb", x"09cc", x"09cc", x"09cc", x"09cc", x"09cd", x"09cd", x"09cd", x"09cd", x"09ce", x"09ce", x"09ce", x"09ce", x"09ce", x"09cf", x"09cf", x"09cf", x"09cf", x"09d0", x"09d0", x"09d0", x"09d0", x"09d1", x"09d1", x"09d1", x"09d1", x"09d2", x"09d2", x"09d2", x"09d2", x"09d2", x"09d3", x"09d3", x"09d3", x"09d3", x"09d4", x"09d4", x"09d4", x"09d4", x"09d5", x"09d5", x"09d5", x"09d5", x"09d6", x"09d6", x"09d6", x"09d6", x"09d7", x"09d7", x"09d7", x"09d7", x"09d7", x"09d8", x"09d8", x"09d8", x"09d8", x"09d9", x"09d9", x"09d9", x"09d9", x"09da", x"09da", x"09da", x"09da", x"09db", x"09db", x"09db", x"09db", x"09db", x"09dc", x"09dc", x"09dc", x"09dc", x"09dd", x"09dd", x"09dd", x"09dd", x"09de", x"09de", x"09de", x"09de", x"09df", x"09df", x"09df", x"09df", x"09e0", x"09e0", x"09e0", x"09e0", x"09e0", x"09e1", x"09e1", x"09e1", x"09e1", x"09e2", x"09e2", x"09e2", x"09e2", x"09e3", x"09e3", x"09e3", x"09e3", x"09e4", x"09e4", x"09e4", x"09e4", x"09e4", x"09e5", x"09e5", x"09e5", x"09e5", x"09e6", x"09e6", x"09e6", x"09e6", x"09e7", x"09e7", x"09e7", x"09e7", x"09e8", x"09e8", x"09e8", x"09e8", x"09e8", x"09e9", x"09e9", x"09e9", x"09e9", x"09ea", x"09ea", x"09ea", x"09ea", x"09eb", x"09eb", x"09eb", x"09eb", x"09ec", x"09ec", x"09ec", x"09ec", x"09ec", x"09ed", x"09ed", x"09ed", x"09ed", x"09ee", x"09ee", x"09ee", x"09ee", x"09ef", x"09ef", x"09ef", x"09ef", x"09f0", x"09f0", x"09f0", x"09f0", x"09f0", x"09f1", x"09f1", x"09f1", x"09f1", x"09f2", x"09f2", x"09f2", x"09f2", x"09f3", x"09f3", x"09f3", x"09f3", x"09f4", x"09f4", x"09f4", x"09f4", x"09f4", x"09f5", x"09f5", x"09f5", x"09f5", x"09f6", x"09f6", x"09f6", x"09f6", x"09f7", x"09f7", x"09f7", x"09f7", x"09f8", x"09f8", x"09f8", x"09f8", x"09f8", x"09f9", x"09f9", x"09f9", x"09f9", x"09fa", x"09fa", x"09fa", x"09fa", x"09fb", x"09fb", x"09fb", x"09fb", x"09fc", x"09fc", x"09fc", x"09fc", x"09fc", x"09fd", x"09fd", x"09fd", x"09fd", x"09fe", x"09fe", x"09fe", x"09fe", x"09ff", x"09ff", x"09ff", x"09ff", x"09ff", x"0a00", x"0a00", x"0a00", x"0a00", x"0a01", x"0a01", x"0a01", x"0a01", x"0a02", x"0a02", x"0a02", x"0a02", x"0a03", x"0a03", x"0a03", x"0a03", x"0a03", x"0a04", x"0a04", x"0a04", x"0a04", x"0a05", x"0a05", x"0a05", x"0a05", x"0a06", x"0a06", x"0a06", x"0a06", x"0a07", x"0a07", x"0a07", x"0a07", x"0a07", x"0a08", x"0a08", x"0a08", x"0a08", x"0a09", x"0a09", x"0a09", x"0a09", x"0a0a", x"0a0a", x"0a0a", x"0a0a", x"0a0a", x"0a0b", x"0a0b", x"0a0b", x"0a0b", x"0a0c", x"0a0c", x"0a0c", x"0a0c", x"0a0d", x"0a0d", x"0a0d", x"0a0d", x"0a0e", x"0a0e", x"0a0e", x"0a0e", x"0a0e", x"0a0f", x"0a0f", x"0a0f", x"0a0f", x"0a10", x"0a10", x"0a10", x"0a10", x"0a11", x"0a11", x"0a11", x"0a11", x"0a11", x"0a12", x"0a12", x"0a12", x"0a12", x"0a13", x"0a13", x"0a13", x"0a13", x"0a14", x"0a14", x"0a14", x"0a14", x"0a15", x"0a15", x"0a15", x"0a15", x"0a15", x"0a16", x"0a16", x"0a16", x"0a16", x"0a17", x"0a17", x"0a17", x"0a17", x"0a18", x"0a18", x"0a18", x"0a18", x"0a18", x"0a19", x"0a19", x"0a19", x"0a19", x"0a1a", x"0a1a", x"0a1a", x"0a1a", x"0a1b", x"0a1b", x"0a1b", x"0a1b", x"0a1c", x"0a1c", x"0a1c", x"0a1c", x"0a1c", x"0a1d", x"0a1d", x"0a1d", x"0a1d", x"0a1e", x"0a1e", x"0a1e", x"0a1e", x"0a1f", x"0a1f", x"0a1f", x"0a1f", x"0a1f", x"0a20", x"0a20", x"0a20", x"0a20", x"0a21", x"0a21", x"0a21", x"0a21", x"0a22", x"0a22", x"0a22", x"0a22", x"0a22", x"0a23", x"0a23", x"0a23", x"0a23", x"0a24", x"0a24", x"0a24", x"0a24", x"0a25", x"0a25", x"0a25", x"0a25", x"0a25", x"0a26", x"0a26", x"0a26", x"0a26", x"0a27", x"0a27", x"0a27", x"0a27", x"0a28", x"0a28", x"0a28", x"0a28", x"0a29", x"0a29", x"0a29", x"0a29", x"0a29", x"0a2a", x"0a2a", x"0a2a", x"0a2a", x"0a2b", x"0a2b", x"0a2b", x"0a2b", x"0a2c", x"0a2c", x"0a2c", x"0a2c", x"0a2c", x"0a2d", x"0a2d", x"0a2d", x"0a2d", x"0a2e", x"0a2e", x"0a2e", x"0a2e", x"0a2f", x"0a2f", x"0a2f", x"0a2f", x"0a2f", x"0a30", x"0a30", x"0a30", x"0a30", x"0a31", x"0a31", x"0a31", x"0a31", x"0a32", x"0a32", x"0a32", x"0a32", x"0a32", x"0a33", x"0a33", x"0a33", x"0a33", x"0a34", x"0a34", x"0a34", x"0a34", x"0a35", x"0a35", x"0a35", x"0a35", x"0a35", x"0a36", x"0a36", x"0a36", x"0a36", x"0a37", x"0a37", x"0a37", x"0a37", x"0a38", x"0a38", x"0a38", x"0a38", x"0a38", x"0a39", x"0a39", x"0a39", x"0a39", x"0a3a", x"0a3a", x"0a3a", x"0a3a", x"0a3b", x"0a3b", x"0a3b", x"0a3b", x"0a3b", x"0a3c", x"0a3c", x"0a3c", x"0a3c", x"0a3d", x"0a3d", x"0a3d", x"0a3d", x"0a3e", x"0a3e", x"0a3e", x"0a3e", x"0a3e", x"0a3f", x"0a3f", x"0a3f", x"0a3f", x"0a40", x"0a40", x"0a40", x"0a40", x"0a41", x"0a41", x"0a41", x"0a41", x"0a41", x"0a42", x"0a42", x"0a42", x"0a42", x"0a43", x"0a43", x"0a43", x"0a43", x"0a44", x"0a44", x"0a44", x"0a44", x"0a44", x"0a45", x"0a45", x"0a45", x"0a45", x"0a46", x"0a46", x"0a46", x"0a46", x"0a46", x"0a47", x"0a47", x"0a47", x"0a47", x"0a48", x"0a48", x"0a48", x"0a48", x"0a49", x"0a49", x"0a49", x"0a49", x"0a49", x"0a4a", x"0a4a", x"0a4a", x"0a4a", x"0a4b", x"0a4b", x"0a4b", x"0a4b", x"0a4c", x"0a4c", x"0a4c", x"0a4c", x"0a4c", x"0a4d", x"0a4d", x"0a4d", x"0a4d", x"0a4e", x"0a4e", x"0a4e", x"0a4e", x"0a4f", x"0a4f", x"0a4f", x"0a4f", x"0a4f", x"0a50", x"0a50", x"0a50", x"0a50", x"0a51", x"0a51", x"0a51", x"0a51", x"0a51", x"0a52", x"0a52", x"0a52", x"0a52", x"0a53", x"0a53", x"0a53", x"0a53", x"0a54", x"0a54", x"0a54", x"0a54", x"0a54", x"0a55", x"0a55", x"0a55", x"0a55", x"0a56", x"0a56", x"0a56", x"0a56", x"0a57", x"0a57", x"0a57", x"0a57", x"0a57", x"0a58", x"0a58", x"0a58", x"0a58", x"0a59", x"0a59", x"0a59", x"0a59", x"0a59", x"0a5a", x"0a5a", x"0a5a", x"0a5a", x"0a5b", x"0a5b", x"0a5b", x"0a5b", x"0a5c", x"0a5c", x"0a5c", x"0a5c", x"0a5c", x"0a5d", x"0a5d", x"0a5d", x"0a5d", x"0a5e", x"0a5e", x"0a5e", x"0a5e", x"0a5f", x"0a5f", x"0a5f", x"0a5f", x"0a5f", x"0a60", x"0a60", x"0a60", x"0a60", x"0a61", x"0a61", x"0a61", x"0a61", x"0a61", x"0a62", x"0a62", x"0a62", x"0a62", x"0a63", x"0a63", x"0a63", x"0a63", x"0a64", x"0a64", x"0a64", x"0a64", x"0a64", x"0a65", x"0a65", x"0a65", x"0a65", x"0a66", x"0a66", x"0a66", x"0a66", x"0a66", x"0a67", x"0a67", x"0a67", x"0a67", x"0a68", x"0a68", x"0a68", x"0a68", x"0a69", x"0a69", x"0a69", x"0a69", x"0a69", x"0a6a", x"0a6a", x"0a6a", x"0a6a", x"0a6b", x"0a6b", x"0a6b", x"0a6b", x"0a6b", x"0a6c", x"0a6c", x"0a6c", x"0a6c", x"0a6d", x"0a6d", x"0a6d", x"0a6d", x"0a6e", x"0a6e", x"0a6e", x"0a6e", x"0a6e", x"0a6f", x"0a6f", x"0a6f", x"0a6f", x"0a70", x"0a70", x"0a70", x"0a70", x"0a70", x"0a71", x"0a71", x"0a71", x"0a71", x"0a72", x"0a72", x"0a72", x"0a72", x"0a73", x"0a73", x"0a73", x"0a73", x"0a73", x"0a74", x"0a74", x"0a74", x"0a74", x"0a75", x"0a75", x"0a75", x"0a75", x"0a75", x"0a76", x"0a76", x"0a76", x"0a76", x"0a77", x"0a77", x"0a77", x"0a77", x"0a77", x"0a78", x"0a78", x"0a78", x"0a78", x"0a79", x"0a79", x"0a79", x"0a79", x"0a7a", x"0a7a", x"0a7a", x"0a7a", x"0a7a", x"0a7b", x"0a7b", x"0a7b", x"0a7b", x"0a7c", x"0a7c", x"0a7c", x"0a7c", x"0a7c", x"0a7d", x"0a7d", x"0a7d", x"0a7d", x"0a7e", x"0a7e", x"0a7e", x"0a7e", x"0a7e", x"0a7f", x"0a7f", x"0a7f", x"0a7f", x"0a80", x"0a80", x"0a80", x"0a80", x"0a81", x"0a81", x"0a81", x"0a81", x"0a81", x"0a82", x"0a82", x"0a82", x"0a82", x"0a83", x"0a83", x"0a83", x"0a83", x"0a83", x"0a84", x"0a84", x"0a84", x"0a84", x"0a85", x"0a85", x"0a85", x"0a85", x"0a85", x"0a86", x"0a86", x"0a86", x"0a86", x"0a87", x"0a87", x"0a87", x"0a87", x"0a87", x"0a88", x"0a88", x"0a88", x"0a88", x"0a89", x"0a89", x"0a89", x"0a89", x"0a8a", x"0a8a", x"0a8a", x"0a8a", x"0a8a", x"0a8b", x"0a8b", x"0a8b", x"0a8b", x"0a8c", x"0a8c", x"0a8c", x"0a8c", x"0a8c", x"0a8d", x"0a8d", x"0a8d", x"0a8d", x"0a8e", x"0a8e", x"0a8e", x"0a8e", x"0a8e", x"0a8f", x"0a8f", x"0a8f", x"0a8f", x"0a90", x"0a90", x"0a90", x"0a90", x"0a90", x"0a91", x"0a91", x"0a91", x"0a91", x"0a92", x"0a92", x"0a92", x"0a92", x"0a92", x"0a93", x"0a93", x"0a93", x"0a93", x"0a94", x"0a94", x"0a94", x"0a94", x"0a95", x"0a95", x"0a95", x"0a95", x"0a95", x"0a96", x"0a96", x"0a96", x"0a96", x"0a97", x"0a97", x"0a97", x"0a97", x"0a97", x"0a98", x"0a98", x"0a98", x"0a98", x"0a99", x"0a99", x"0a99", x"0a99", x"0a99", x"0a9a", x"0a9a", x"0a9a", x"0a9a", x"0a9b", x"0a9b", x"0a9b", x"0a9b", x"0a9b", x"0a9c", x"0a9c", x"0a9c", x"0a9c", x"0a9d", x"0a9d", x"0a9d", x"0a9d", x"0a9d", x"0a9e", x"0a9e", x"0a9e", x"0a9e", x"0a9f", x"0a9f", x"0a9f", x"0a9f", x"0a9f", x"0aa0", x"0aa0", x"0aa0", x"0aa0", x"0aa1", x"0aa1", x"0aa1", x"0aa1", x"0aa1", x"0aa2", x"0aa2", x"0aa2", x"0aa2", x"0aa3", x"0aa3", x"0aa3", x"0aa3", x"0aa3", x"0aa4", x"0aa4", x"0aa4", x"0aa4", x"0aa5", x"0aa5", x"0aa5", x"0aa5", x"0aa5", x"0aa6", x"0aa6", x"0aa6", x"0aa6", x"0aa7", x"0aa7", x"0aa7", x"0aa7", x"0aa7", x"0aa8", x"0aa8", x"0aa8", x"0aa8", x"0aa9", x"0aa9", x"0aa9", x"0aa9", x"0aa9", x"0aaa", x"0aaa", x"0aaa", x"0aaa", x"0aab", x"0aab", x"0aab", x"0aab", x"0aab", x"0aac", x"0aac", x"0aac", x"0aac", x"0aad", x"0aad", x"0aad", x"0aad", x"0aad", x"0aae", x"0aae", x"0aae", x"0aae", x"0aaf", x"0aaf", x"0aaf", x"0aaf", x"0aaf", x"0ab0", x"0ab0", x"0ab0", x"0ab0", x"0ab1", x"0ab1", x"0ab1", x"0ab1", x"0ab1", x"0ab2", x"0ab2", x"0ab2", x"0ab2", x"0ab3", x"0ab3", x"0ab3", x"0ab3", x"0ab3", x"0ab4", x"0ab4", x"0ab4", x"0ab4", x"0ab5", x"0ab5", x"0ab5", x"0ab5", x"0ab5", x"0ab6", x"0ab6", x"0ab6", x"0ab6", x"0ab7", x"0ab7", x"0ab7", x"0ab7", x"0ab7", x"0ab8", x"0ab8", x"0ab8", x"0ab8", x"0ab9", x"0ab9", x"0ab9", x"0ab9", x"0ab9", x"0aba", x"0aba", x"0aba", x"0aba", x"0abb", x"0abb", x"0abb", x"0abb", x"0abb", x"0abc", x"0abc", x"0abc", x"0abc", x"0abd", x"0abd", x"0abd", x"0abd", x"0abd", x"0abe", x"0abe", x"0abe", x"0abe", x"0abe", x"0abf", x"0abf", x"0abf", x"0abf", x"0ac0", x"0ac0", x"0ac0", x"0ac0", x"0ac0", x"0ac1", x"0ac1", x"0ac1", x"0ac1", x"0ac2", x"0ac2", x"0ac2", x"0ac2", x"0ac2", x"0ac3", x"0ac3", x"0ac3", x"0ac3", x"0ac4", x"0ac4", x"0ac4", x"0ac4", x"0ac4", x"0ac5", x"0ac5", x"0ac5", x"0ac5", x"0ac6", x"0ac6", x"0ac6", x"0ac6", x"0ac6", x"0ac7", x"0ac7", x"0ac7", x"0ac7", x"0ac8", x"0ac8", x"0ac8", x"0ac8", x"0ac8", x"0ac9", x"0ac9", x"0ac9", x"0ac9", x"0ac9", x"0aca", x"0aca", x"0aca", x"0aca", x"0acb", x"0acb", x"0acb", x"0acb", x"0acb", x"0acc", x"0acc", x"0acc", x"0acc", x"0acd", x"0acd", x"0acd", x"0acd", x"0acd", x"0ace", x"0ace", x"0ace", x"0ace", x"0acf", x"0acf", x"0acf", x"0acf", x"0acf", x"0ad0", x"0ad0", x"0ad0", x"0ad0", x"0ad1", x"0ad1", x"0ad1", x"0ad1", x"0ad1", x"0ad2", x"0ad2", x"0ad2", x"0ad2", x"0ad2", x"0ad3", x"0ad3", x"0ad3", x"0ad3", x"0ad4", x"0ad4", x"0ad4", x"0ad4", x"0ad4", x"0ad5", x"0ad5", x"0ad5", x"0ad5", x"0ad6", x"0ad6", x"0ad6", x"0ad6", x"0ad6", x"0ad7", x"0ad7", x"0ad7", x"0ad7", x"0ad8", x"0ad8", x"0ad8", x"0ad8", x"0ad8", x"0ad9", x"0ad9", x"0ad9", x"0ad9", x"0ad9", x"0ada", x"0ada", x"0ada", x"0ada", x"0adb", x"0adb", x"0adb", x"0adb", x"0adb", x"0adc", x"0adc", x"0adc", x"0adc", x"0add", x"0add", x"0add", x"0add", x"0add", x"0ade", x"0ade", x"0ade", x"0ade", x"0ade", x"0adf", x"0adf", x"0adf", x"0adf", x"0ae0", x"0ae0", x"0ae0", x"0ae0", x"0ae0", x"0ae1", x"0ae1", x"0ae1", x"0ae1", x"0ae2", x"0ae2", x"0ae2", x"0ae2", x"0ae2", x"0ae3", x"0ae3", x"0ae3", x"0ae3", x"0ae3", x"0ae4", x"0ae4", x"0ae4", x"0ae4", x"0ae5", x"0ae5", x"0ae5", x"0ae5", x"0ae5", x"0ae6", x"0ae6", x"0ae6", x"0ae6", x"0ae7", x"0ae7", x"0ae7", x"0ae7", x"0ae7", x"0ae8", x"0ae8", x"0ae8", x"0ae8", x"0ae8", x"0ae9", x"0ae9", x"0ae9", x"0ae9", x"0aea", x"0aea", x"0aea", x"0aea", x"0aea", x"0aeb", x"0aeb", x"0aeb", x"0aeb", x"0aec", x"0aec", x"0aec", x"0aec", x"0aec", x"0aed", x"0aed", x"0aed", x"0aed", x"0aed", x"0aee", x"0aee", x"0aee", x"0aee", x"0aef", x"0aef", x"0aef", x"0aef", x"0aef", x"0af0", x"0af0", x"0af0", x"0af0", x"0af0", x"0af1", x"0af1", x"0af1", x"0af1", x"0af2", x"0af2", x"0af2", x"0af2", x"0af2", x"0af3", x"0af3", x"0af3", x"0af3", x"0af4", x"0af4", x"0af4", x"0af4", x"0af4", x"0af5", x"0af5", x"0af5", x"0af5", x"0af5", x"0af6", x"0af6", x"0af6", x"0af6", x"0af7", x"0af7", x"0af7", x"0af7", x"0af7", x"0af8", x"0af8", x"0af8", x"0af8", x"0af8", x"0af9", x"0af9", x"0af9", x"0af9", x"0afa", x"0afa", x"0afa", x"0afa", x"0afa", x"0afb", x"0afb", x"0afb", x"0afb", x"0afb", x"0afc", x"0afc", x"0afc", x"0afc", x"0afd", x"0afd", x"0afd", x"0afd", x"0afd", x"0afe", x"0afe", x"0afe", x"0afe", x"0afe", x"0aff", x"0aff", x"0aff", x"0aff", x"0b00", x"0b00", x"0b00", x"0b00", x"0b00", x"0b01", x"0b01", x"0b01", x"0b01", x"0b01", x"0b02", x"0b02", x"0b02", x"0b02", x"0b03", x"0b03", x"0b03", x"0b03", x"0b03", x"0b04", x"0b04", x"0b04", x"0b04", x"0b04", x"0b05", x"0b05", x"0b05", x"0b05", x"0b06", x"0b06", x"0b06", x"0b06", x"0b06", x"0b07", x"0b07", x"0b07", x"0b07", x"0b07", x"0b08", x"0b08", x"0b08", x"0b08", x"0b09", x"0b09", x"0b09", x"0b09", x"0b09", x"0b0a", x"0b0a", x"0b0a", x"0b0a", x"0b0a", x"0b0b", x"0b0b", x"0b0b", x"0b0b", x"0b0c", x"0b0c", x"0b0c", x"0b0c", x"0b0c", x"0b0d", x"0b0d", x"0b0d", x"0b0d", x"0b0d", x"0b0e", x"0b0e", x"0b0e", x"0b0e", x"0b0f", x"0b0f", x"0b0f", x"0b0f", x"0b0f", x"0b10", x"0b10", x"0b10", x"0b10", x"0b10", x"0b11", x"0b11", x"0b11", x"0b11", x"0b12", x"0b12", x"0b12", x"0b12", x"0b12", x"0b13", x"0b13", x"0b13", x"0b13", x"0b13", x"0b14", x"0b14", x"0b14", x"0b14", x"0b15", x"0b15", x"0b15", x"0b15", x"0b15", x"0b16", x"0b16", x"0b16", x"0b16", x"0b16", x"0b17", x"0b17", x"0b17", x"0b17", x"0b17", x"0b18", x"0b18", x"0b18", x"0b18", x"0b19", x"0b19", x"0b19", x"0b19", x"0b19", x"0b1a", x"0b1a", x"0b1a", x"0b1a", x"0b1a", x"0b1b", x"0b1b", x"0b1b", x"0b1b", x"0b1c", x"0b1c", x"0b1c", x"0b1c", x"0b1c", x"0b1d", x"0b1d", x"0b1d", x"0b1d", x"0b1d", x"0b1e", x"0b1e", x"0b1e", x"0b1e", x"0b1e", x"0b1f", x"0b1f", x"0b1f", x"0b1f", x"0b20", x"0b20", x"0b20", x"0b20", x"0b20", x"0b21", x"0b21", x"0b21", x"0b21", x"0b21", x"0b22", x"0b22", x"0b22", x"0b22", x"0b23", x"0b23", x"0b23", x"0b23", x"0b23", x"0b24", x"0b24", x"0b24", x"0b24", x"0b24", x"0b25", x"0b25", x"0b25", x"0b25", x"0b25", x"0b26", x"0b26", x"0b26", x"0b26", x"0b27", x"0b27", x"0b27", x"0b27", x"0b27", x"0b28", x"0b28", x"0b28", x"0b28", x"0b28", x"0b29", x"0b29", x"0b29", x"0b29", x"0b29", x"0b2a", x"0b2a", x"0b2a", x"0b2a", x"0b2b", x"0b2b", x"0b2b", x"0b2b", x"0b2b", x"0b2c", x"0b2c", x"0b2c", x"0b2c", x"0b2c", x"0b2d", x"0b2d", x"0b2d", x"0b2d", x"0b2d", x"0b2e", x"0b2e", x"0b2e", x"0b2e", x"0b2f", x"0b2f", x"0b2f", x"0b2f", x"0b2f", x"0b30", x"0b30", x"0b30", x"0b30", x"0b30", x"0b31", x"0b31", x"0b31", x"0b31", x"0b31", x"0b32", x"0b32", x"0b32", x"0b32", x"0b33", x"0b33", x"0b33", x"0b33", x"0b33", x"0b34", x"0b34", x"0b34", x"0b34", x"0b34", x"0b35", x"0b35", x"0b35", x"0b35", x"0b35", x"0b36", x"0b36", x"0b36", x"0b36", x"0b37", x"0b37", x"0b37", x"0b37", x"0b37", x"0b38", x"0b38", x"0b38", x"0b38", x"0b38", x"0b39", x"0b39", x"0b39", x"0b39", x"0b39", x"0b3a", x"0b3a", x"0b3a", x"0b3a", x"0b3a", x"0b3b", x"0b3b", x"0b3b", x"0b3b", x"0b3c", x"0b3c", x"0b3c", x"0b3c", x"0b3c", x"0b3d", x"0b3d", x"0b3d", x"0b3d", x"0b3d", x"0b3e", x"0b3e", x"0b3e", x"0b3e", x"0b3e", x"0b3f", x"0b3f", x"0b3f", x"0b3f", x"0b3f", x"0b40", x"0b40", x"0b40", x"0b40", x"0b41", x"0b41", x"0b41", x"0b41", x"0b41", x"0b42", x"0b42", x"0b42", x"0b42", x"0b42", x"0b43", x"0b43", x"0b43", x"0b43", x"0b43", x"0b44", x"0b44", x"0b44", x"0b44", x"0b44", x"0b45", x"0b45", x"0b45", x"0b45", x"0b46", x"0b46", x"0b46", x"0b46", x"0b46", x"0b47", x"0b47", x"0b47", x"0b47", x"0b47", x"0b48", x"0b48", x"0b48", x"0b48", x"0b48", x"0b49", x"0b49", x"0b49", x"0b49", x"0b49", x"0b4a", x"0b4a", x"0b4a", x"0b4a", x"0b4b", x"0b4b", x"0b4b", x"0b4b", x"0b4b", x"0b4c", x"0b4c", x"0b4c", x"0b4c", x"0b4c", x"0b4d", x"0b4d", x"0b4d", x"0b4d", x"0b4d", x"0b4e", x"0b4e", x"0b4e", x"0b4e", x"0b4e", x"0b4f", x"0b4f", x"0b4f", x"0b4f", x"0b4f", x"0b50", x"0b50", x"0b50", x"0b50", x"0b51", x"0b51", x"0b51", x"0b51", x"0b51", x"0b52", x"0b52", x"0b52", x"0b52", x"0b52", x"0b53", x"0b53", x"0b53", x"0b53", x"0b53", x"0b54", x"0b54", x"0b54", x"0b54", x"0b54", x"0b55", x"0b55", x"0b55", x"0b55", x"0b55", x"0b56", x"0b56", x"0b56", x"0b56", x"0b57", x"0b57", x"0b57", x"0b57", x"0b57", x"0b58", x"0b58", x"0b58", x"0b58", x"0b58", x"0b59", x"0b59", x"0b59", x"0b59", x"0b59", x"0b5a", x"0b5a", x"0b5a", x"0b5a", x"0b5a", x"0b5b", x"0b5b", x"0b5b", x"0b5b", x"0b5b", x"0b5c", x"0b5c", x"0b5c", x"0b5c", x"0b5c", x"0b5d", x"0b5d", x"0b5d", x"0b5d", x"0b5e", x"0b5e", x"0b5e", x"0b5e", x"0b5e", x"0b5f", x"0b5f", x"0b5f", x"0b5f", x"0b5f", x"0b60", x"0b60", x"0b60", x"0b60", x"0b60", x"0b61", x"0b61", x"0b61", x"0b61", x"0b61", x"0b62", x"0b62", x"0b62", x"0b62", x"0b62", x"0b63", x"0b63", x"0b63", x"0b63", x"0b63", x"0b64", x"0b64", x"0b64", x"0b64", x"0b65", x"0b65", x"0b65", x"0b65", x"0b65", x"0b66", x"0b66", x"0b66", x"0b66", x"0b66", x"0b67", x"0b67", x"0b67", x"0b67", x"0b67", x"0b68", x"0b68", x"0b68", x"0b68", x"0b68", x"0b69", x"0b69", x"0b69", x"0b69", x"0b69", x"0b6a", x"0b6a", x"0b6a", x"0b6a", x"0b6a", x"0b6b", x"0b6b", x"0b6b", x"0b6b", x"0b6b", x"0b6c", x"0b6c", x"0b6c", x"0b6c", x"0b6c", x"0b6d", x"0b6d", x"0b6d", x"0b6d", x"0b6d", x"0b6e", x"0b6e", x"0b6e", x"0b6e", x"0b6f", x"0b6f", x"0b6f", x"0b6f", x"0b6f", x"0b70", x"0b70", x"0b70", x"0b70", x"0b70", x"0b71", x"0b71", x"0b71", x"0b71", x"0b71", x"0b72", x"0b72", x"0b72", x"0b72", x"0b72", x"0b73", x"0b73", x"0b73", x"0b73", x"0b73", x"0b74", x"0b74", x"0b74", x"0b74", x"0b74", x"0b75", x"0b75", x"0b75", x"0b75", x"0b75", x"0b76", x"0b76", x"0b76", x"0b76", x"0b76", x"0b77", x"0b77", x"0b77", x"0b77", x"0b77", x"0b78", x"0b78", x"0b78", x"0b78", x"0b78", x"0b79", x"0b79", x"0b79", x"0b79", x"0b79", x"0b7a", x"0b7a", x"0b7a", x"0b7a", x"0b7b", x"0b7b", x"0b7b", x"0b7b", x"0b7b", x"0b7c", x"0b7c", x"0b7c", x"0b7c", x"0b7c", x"0b7d", x"0b7d", x"0b7d", x"0b7d", x"0b7d", x"0b7e", x"0b7e", x"0b7e", x"0b7e", x"0b7e", x"0b7f", x"0b7f", x"0b7f", x"0b7f", x"0b7f", x"0b80", x"0b80", x"0b80", x"0b80", x"0b80", x"0b81", x"0b81", x"0b81", x"0b81", x"0b81", x"0b82", x"0b82", x"0b82", x"0b82", x"0b82", x"0b83", x"0b83", x"0b83", x"0b83", x"0b83", x"0b84", x"0b84", x"0b84", x"0b84", x"0b84", x"0b85", x"0b85", x"0b85", x"0b85", x"0b85", x"0b86", x"0b86", x"0b86", x"0b86", x"0b86", x"0b87", x"0b87", x"0b87", x"0b87", x"0b87", x"0b88", x"0b88", x"0b88", x"0b88", x"0b88", x"0b89", x"0b89", x"0b89", x"0b89", x"0b89", x"0b8a", x"0b8a", x"0b8a", x"0b8a", x"0b8a", x"0b8b", x"0b8b", x"0b8b", x"0b8b", x"0b8b", x"0b8c", x"0b8c", x"0b8c", x"0b8c", x"0b8c", x"0b8d", x"0b8d", x"0b8d", x"0b8d", x"0b8d", x"0b8e", x"0b8e", x"0b8e", x"0b8e", x"0b8e", x"0b8f", x"0b8f", x"0b8f", x"0b8f", x"0b8f", x"0b90", x"0b90", x"0b90", x"0b90", x"0b90", x"0b91", x"0b91", x"0b91", x"0b91", x"0b91", x"0b92", x"0b92", x"0b92", x"0b92", x"0b92", x"0b93", x"0b93", x"0b93", x"0b93", x"0b93", x"0b94", x"0b94", x"0b94", x"0b94", x"0b94", x"0b95", x"0b95", x"0b95", x"0b95", x"0b95", x"0b96", x"0b96", x"0b96", x"0b96", x"0b96", x"0b97", x"0b97", x"0b97", x"0b97", x"0b97", x"0b98", x"0b98", x"0b98", x"0b98", x"0b98", x"0b99", x"0b99", x"0b99", x"0b99", x"0b99", x"0b9a", x"0b9a", x"0b9a", x"0b9a", x"0b9a", x"0b9b", x"0b9b", x"0b9b", x"0b9b", x"0b9b", x"0b9c", x"0b9c", x"0b9c", x"0b9c", x"0b9c", x"0b9d", x"0b9d", x"0b9d", x"0b9d", x"0b9d", x"0b9e", x"0b9e", x"0b9e", x"0b9e", x"0b9e", x"0b9f", x"0b9f", x"0b9f", x"0b9f", x"0b9f", x"0ba0", x"0ba0", x"0ba0", x"0ba0", x"0ba0", x"0ba1", x"0ba1", x"0ba1", x"0ba1", x"0ba1", x"0ba2", x"0ba2", x"0ba2", x"0ba2", x"0ba2", x"0ba3", x"0ba3", x"0ba3", x"0ba3", x"0ba3", x"0ba4", x"0ba4", x"0ba4", x"0ba4", x"0ba4", x"0ba5", x"0ba5", x"0ba5", x"0ba5", x"0ba5", x"0ba6", x"0ba6", x"0ba6", x"0ba6", x"0ba6", x"0ba7", x"0ba7", x"0ba7", x"0ba7", x"0ba7", x"0ba8", x"0ba8", x"0ba8", x"0ba8", x"0ba8", x"0ba9", x"0ba9", x"0ba9", x"0ba9", x"0ba9", x"0baa", x"0baa", x"0baa", x"0baa", x"0baa", x"0baa", x"0bab", x"0bab", x"0bab", x"0bab", x"0bab", x"0bac", x"0bac", x"0bac", x"0bac", x"0bac", x"0bad", x"0bad", x"0bad", x"0bad", x"0bad", x"0bae", x"0bae", x"0bae", x"0bae", x"0bae", x"0baf", x"0baf", x"0baf", x"0baf", x"0baf", x"0bb0", x"0bb0", x"0bb0", x"0bb0", x"0bb0", x"0bb1", x"0bb1", x"0bb1", x"0bb1", x"0bb1", x"0bb2", x"0bb2", x"0bb2", x"0bb2", x"0bb2", x"0bb3", x"0bb3", x"0bb3", x"0bb3", x"0bb3", x"0bb4", x"0bb4", x"0bb4", x"0bb4", x"0bb4", x"0bb5", x"0bb5", x"0bb5", x"0bb5", x"0bb5", x"0bb6", x"0bb6", x"0bb6", x"0bb6", x"0bb6", x"0bb6", x"0bb7", x"0bb7", x"0bb7", x"0bb7", x"0bb7", x"0bb8", x"0bb8", x"0bb8", x"0bb8", x"0bb8", x"0bb9", x"0bb9", x"0bb9", x"0bb9", x"0bb9", x"0bba", x"0bba", x"0bba", x"0bba", x"0bba", x"0bbb", x"0bbb", x"0bbb", x"0bbb", x"0bbb", x"0bbc", x"0bbc", x"0bbc", x"0bbc", x"0bbc", x"0bbd", x"0bbd", x"0bbd", x"0bbd", x"0bbd", x"0bbe", x"0bbe", x"0bbe", x"0bbe", x"0bbe", x"0bbe", x"0bbf", x"0bbf", x"0bbf", x"0bbf", x"0bbf", x"0bc0", x"0bc0", x"0bc0", x"0bc0", x"0bc0", x"0bc1", x"0bc1", x"0bc1", x"0bc1", x"0bc1", x"0bc2", x"0bc2", x"0bc2", x"0bc2", x"0bc2", x"0bc3", x"0bc3", x"0bc3", x"0bc3", x"0bc3", x"0bc4", x"0bc4", x"0bc4", x"0bc4", x"0bc4", x"0bc5", x"0bc5", x"0bc5", x"0bc5", x"0bc5", x"0bc6", x"0bc6", x"0bc6", x"0bc6", x"0bc6", x"0bc6", x"0bc7", x"0bc7", x"0bc7", x"0bc7", x"0bc7", x"0bc8", x"0bc8", x"0bc8", x"0bc8", x"0bc8", x"0bc9", x"0bc9", x"0bc9", x"0bc9", x"0bc9", x"0bca", x"0bca", x"0bca", x"0bca", x"0bca", x"0bcb", x"0bcb", x"0bcb", x"0bcb", x"0bcb", x"0bcc", x"0bcc", x"0bcc", x"0bcc", x"0bcc", x"0bcc", x"0bcd", x"0bcd", x"0bcd", x"0bcd", x"0bcd", x"0bce", x"0bce", x"0bce", x"0bce", x"0bce", x"0bcf", x"0bcf", x"0bcf", x"0bcf", x"0bcf", x"0bd0", x"0bd0", x"0bd0", x"0bd0", x"0bd0", x"0bd1", x"0bd1", x"0bd1", x"0bd1", x"0bd1", x"0bd2", x"0bd2", x"0bd2", x"0bd2", x"0bd2", x"0bd2", x"0bd3", x"0bd3", x"0bd3", x"0bd3", x"0bd3", x"0bd4", x"0bd4", x"0bd4", x"0bd4", x"0bd4", x"0bd5", x"0bd5", x"0bd5", x"0bd5", x"0bd5", x"0bd6", x"0bd6", x"0bd6", x"0bd6", x"0bd6", x"0bd7", x"0bd7", x"0bd7", x"0bd7", x"0bd7", x"0bd7", x"0bd8", x"0bd8", x"0bd8", x"0bd8", x"0bd8", x"0bd9", x"0bd9", x"0bd9", x"0bd9", x"0bd9", x"0bda", x"0bda", x"0bda", x"0bda", x"0bda", x"0bdb", x"0bdb", x"0bdb", x"0bdb", x"0bdb", x"0bdc", x"0bdc", x"0bdc", x"0bdc", x"0bdc", x"0bdc", x"0bdd", x"0bdd", x"0bdd", x"0bdd", x"0bdd", x"0bde", x"0bde", x"0bde", x"0bde", x"0bde", x"0bdf", x"0bdf", x"0bdf", x"0bdf", x"0bdf", x"0be0", x"0be0", x"0be0", x"0be0", x"0be0", x"0be0", x"0be1", x"0be1", x"0be1", x"0be1", x"0be1", x"0be2", x"0be2", x"0be2", x"0be2", x"0be2", x"0be3", x"0be3", x"0be3", x"0be3", x"0be3", x"0be4", x"0be4", x"0be4", x"0be4", x"0be4", x"0be4", x"0be5", x"0be5", x"0be5", x"0be5", x"0be5", x"0be6", x"0be6", x"0be6", x"0be6", x"0be6", x"0be7", x"0be7", x"0be7", x"0be7", x"0be7", x"0be8", x"0be8", x"0be8", x"0be8", x"0be8", x"0be8", x"0be9", x"0be9", x"0be9", x"0be9", x"0be9", x"0bea", x"0bea", x"0bea", x"0bea", x"0bea", x"0beb", x"0beb", x"0beb", x"0beb", x"0beb", x"0bec", x"0bec", x"0bec", x"0bec", x"0bec", x"0bec", x"0bed", x"0bed", x"0bed", x"0bed", x"0bed", x"0bee", x"0bee", x"0bee", x"0bee", x"0bee", x"0bef", x"0bef", x"0bef", x"0bef", x"0bef", x"0bf0", x"0bf0", x"0bf0", x"0bf0", x"0bf0", x"0bf0", x"0bf1", x"0bf1", x"0bf1", x"0bf1", x"0bf1", x"0bf2", x"0bf2", x"0bf2", x"0bf2", x"0bf2", x"0bf3", x"0bf3", x"0bf3", x"0bf3", x"0bf3", x"0bf3", x"0bf4", x"0bf4", x"0bf4", x"0bf4", x"0bf4", x"0bf5", x"0bf5", x"0bf5", x"0bf5", x"0bf5", x"0bf6", x"0bf6", x"0bf6", x"0bf6", x"0bf6", x"0bf6", x"0bf7", x"0bf7", x"0bf7", x"0bf7", x"0bf7", x"0bf8", x"0bf8", x"0bf8", x"0bf8", x"0bf8", x"0bf9", x"0bf9", x"0bf9", x"0bf9", x"0bf9", x"0bfa", x"0bfa", x"0bfa", x"0bfa", x"0bfa", x"0bfa", x"0bfb", x"0bfb", x"0bfb", x"0bfb", x"0bfb", x"0bfc", x"0bfc", x"0bfc", x"0bfc", x"0bfc", x"0bfd", x"0bfd", x"0bfd", x"0bfd", x"0bfd", x"0bfd", x"0bfe", x"0bfe", x"0bfe", x"0bfe", x"0bfe", x"0bff", x"0bff", x"0bff", x"0bff", x"0bff", x"0c00", x"0c00", x"0c00", x"0c00", x"0c00", x"0c00", x"0c01", x"0c01", x"0c01", x"0c01", x"0c01", x"0c02", x"0c02", x"0c02", x"0c02", x"0c02", x"0c03", x"0c03", x"0c03", x"0c03", x"0c03", x"0c03", x"0c04", x"0c04", x"0c04", x"0c04", x"0c04", x"0c05", x"0c05", x"0c05", x"0c05", x"0c05", x"0c05", x"0c06", x"0c06", x"0c06", x"0c06", x"0c06", x"0c07", x"0c07", x"0c07", x"0c07", x"0c07", x"0c08", x"0c08", x"0c08", x"0c08", x"0c08", x"0c08", x"0c09", x"0c09", x"0c09", x"0c09", x"0c09", x"0c0a", x"0c0a", x"0c0a", x"0c0a", x"0c0a", x"0c0b", x"0c0b", x"0c0b", x"0c0b", x"0c0b", x"0c0b", x"0c0c", x"0c0c", x"0c0c", x"0c0c", x"0c0c", x"0c0d", x"0c0d", x"0c0d", x"0c0d", x"0c0d", x"0c0e", x"0c0e", x"0c0e", x"0c0e", x"0c0e", x"0c0e", x"0c0f", x"0c0f", x"0c0f", x"0c0f", x"0c0f", x"0c10", x"0c10", x"0c10", x"0c10", x"0c10", x"0c10", x"0c11", x"0c11", x"0c11", x"0c11", x"0c11", x"0c12", x"0c12", x"0c12", x"0c12", x"0c12", x"0c13", x"0c13", x"0c13", x"0c13", x"0c13", x"0c13", x"0c14", x"0c14", x"0c14", x"0c14", x"0c14", x"0c15", x"0c15", x"0c15", x"0c15", x"0c15", x"0c15", x"0c16", x"0c16", x"0c16", x"0c16", x"0c16", x"0c17", x"0c17", x"0c17", x"0c17", x"0c17", x"0c17", x"0c18", x"0c18", x"0c18", x"0c18", x"0c18", x"0c19", x"0c19", x"0c19", x"0c19", x"0c19", x"0c1a", x"0c1a", x"0c1a", x"0c1a", x"0c1a", x"0c1a", x"0c1b", x"0c1b", x"0c1b", x"0c1b", x"0c1b", x"0c1c", x"0c1c", x"0c1c", x"0c1c", x"0c1c", x"0c1c", x"0c1d", x"0c1d", x"0c1d", x"0c1d", x"0c1d", x"0c1e", x"0c1e", x"0c1e", x"0c1e", x"0c1e", x"0c1e", x"0c1f", x"0c1f", x"0c1f", x"0c1f", x"0c1f", x"0c20", x"0c20", x"0c20", x"0c20", x"0c20", x"0c21", x"0c21", x"0c21", x"0c21", x"0c21", x"0c21", x"0c22", x"0c22", x"0c22", x"0c22", x"0c22", x"0c23", x"0c23", x"0c23", x"0c23", x"0c23", x"0c23", x"0c24", x"0c24", x"0c24", x"0c24", x"0c24", x"0c25", x"0c25", x"0c25", x"0c25", x"0c25", x"0c25", x"0c26", x"0c26", x"0c26", x"0c26", x"0c26", x"0c27", x"0c27", x"0c27", x"0c27", x"0c27", x"0c27", x"0c28", x"0c28", x"0c28", x"0c28", x"0c28", x"0c29", x"0c29", x"0c29", x"0c29", x"0c29", x"0c29", x"0c2a", x"0c2a", x"0c2a", x"0c2a", x"0c2a", x"0c2b", x"0c2b", x"0c2b", x"0c2b", x"0c2b", x"0c2b", x"0c2c", x"0c2c", x"0c2c", x"0c2c", x"0c2c", x"0c2d", x"0c2d", x"0c2d", x"0c2d", x"0c2d", x"0c2d", x"0c2e", x"0c2e", x"0c2e", x"0c2e", x"0c2e", x"0c2f", x"0c2f", x"0c2f", x"0c2f", x"0c2f", x"0c2f", x"0c30", x"0c30", x"0c30", x"0c30", x"0c30", x"0c31", x"0c31", x"0c31", x"0c31", x"0c31", x"0c31", x"0c32", x"0c32", x"0c32", x"0c32", x"0c32", x"0c33", x"0c33", x"0c33", x"0c33", x"0c33", x"0c33", x"0c34", x"0c34", x"0c34", x"0c34", x"0c34", x"0c35", x"0c35", x"0c35", x"0c35", x"0c35", x"0c35", x"0c36", x"0c36", x"0c36", x"0c36", x"0c36", x"0c37", x"0c37", x"0c37", x"0c37", x"0c37", x"0c37", x"0c38", x"0c38", x"0c38", x"0c38", x"0c38", x"0c38", x"0c39", x"0c39", x"0c39", x"0c39", x"0c39", x"0c3a", x"0c3a", x"0c3a", x"0c3a", x"0c3a", x"0c3a", x"0c3b", x"0c3b", x"0c3b", x"0c3b", x"0c3b", x"0c3c", x"0c3c", x"0c3c", x"0c3c", x"0c3c", x"0c3c", x"0c3d", x"0c3d", x"0c3d", x"0c3d", x"0c3d", x"0c3e", x"0c3e", x"0c3e", x"0c3e", x"0c3e", x"0c3e", x"0c3f", x"0c3f", x"0c3f", x"0c3f", x"0c3f", x"0c40", x"0c40", x"0c40", x"0c40", x"0c40", x"0c40", x"0c41", x"0c41", x"0c41", x"0c41", x"0c41", x"0c41", x"0c42", x"0c42", x"0c42", x"0c42", x"0c42", x"0c43", x"0c43", x"0c43", x"0c43", x"0c43", x"0c43", x"0c44", x"0c44", x"0c44", x"0c44", x"0c44", x"0c45", x"0c45", x"0c45", x"0c45", x"0c45", x"0c45", x"0c46", x"0c46", x"0c46", x"0c46", x"0c46", x"0c46", x"0c47", x"0c47", x"0c47", x"0c47", x"0c47", x"0c48", x"0c48", x"0c48", x"0c48", x"0c48", x"0c48", x"0c49", x"0c49", x"0c49", x"0c49", x"0c49", x"0c4a", x"0c4a", x"0c4a", x"0c4a", x"0c4a", x"0c4a", x"0c4b", x"0c4b", x"0c4b", x"0c4b", x"0c4b", x"0c4b", x"0c4c", x"0c4c", x"0c4c", x"0c4c", x"0c4c", x"0c4d", x"0c4d", x"0c4d", x"0c4d", x"0c4d", x"0c4d", x"0c4e", x"0c4e", x"0c4e", x"0c4e", x"0c4e", x"0c4e", x"0c4f", x"0c4f", x"0c4f", x"0c4f", x"0c4f", x"0c50", x"0c50", x"0c50", x"0c50", x"0c50", x"0c50", x"0c51", x"0c51", x"0c51", x"0c51", x"0c51", x"0c51", x"0c52", x"0c52", x"0c52", x"0c52", x"0c52", x"0c53", x"0c53", x"0c53", x"0c53", x"0c53", x"0c53", x"0c54", x"0c54", x"0c54", x"0c54", x"0c54", x"0c54", x"0c55", x"0c55", x"0c55", x"0c55", x"0c55", x"0c56", x"0c56", x"0c56", x"0c56", x"0c56", x"0c56", x"0c57", x"0c57", x"0c57", x"0c57", x"0c57", x"0c57", x"0c58", x"0c58", x"0c58", x"0c58", x"0c58", x"0c59", x"0c59", x"0c59", x"0c59", x"0c59", x"0c59", x"0c5a", x"0c5a", x"0c5a", x"0c5a", x"0c5a", x"0c5a", x"0c5b", x"0c5b", x"0c5b", x"0c5b", x"0c5b", x"0c5c", x"0c5c", x"0c5c", x"0c5c", x"0c5c", x"0c5c", x"0c5d", x"0c5d", x"0c5d", x"0c5d", x"0c5d", x"0c5d", x"0c5e", x"0c5e", x"0c5e", x"0c5e", x"0c5e", x"0c5f", x"0c5f", x"0c5f", x"0c5f", x"0c5f", x"0c5f", x"0c60", x"0c60", x"0c60", x"0c60", x"0c60", x"0c60", x"0c61", x"0c61", x"0c61", x"0c61", x"0c61", x"0c61", x"0c62", x"0c62", x"0c62", x"0c62", x"0c62", x"0c63", x"0c63", x"0c63", x"0c63", x"0c63", x"0c63", x"0c64", x"0c64", x"0c64", x"0c64", x"0c64", x"0c64", x"0c65", x"0c65", x"0c65", x"0c65", x"0c65", x"0c66", x"0c66", x"0c66", x"0c66", x"0c66", x"0c66", x"0c67", x"0c67", x"0c67", x"0c67", x"0c67", x"0c67", x"0c68", x"0c68", x"0c68", x"0c68", x"0c68", x"0c68", x"0c69", x"0c69", x"0c69", x"0c69", x"0c69", x"0c6a", x"0c6a", x"0c6a", x"0c6a", x"0c6a", x"0c6a", x"0c6b", x"0c6b", x"0c6b", x"0c6b", x"0c6b", x"0c6b", x"0c6c", x"0c6c", x"0c6c", x"0c6c", x"0c6c", x"0c6c", x"0c6d", x"0c6d", x"0c6d", x"0c6d", x"0c6d", x"0c6e", x"0c6e", x"0c6e", x"0c6e", x"0c6e", x"0c6e", x"0c6f", x"0c6f", x"0c6f", x"0c6f", x"0c6f", x"0c6f", x"0c70", x"0c70", x"0c70", x"0c70", x"0c70", x"0c70", x"0c71", x"0c71", x"0c71", x"0c71", x"0c71", x"0c71", x"0c72", x"0c72", x"0c72", x"0c72", x"0c72", x"0c73", x"0c73", x"0c73", x"0c73", x"0c73", x"0c73", x"0c74", x"0c74", x"0c74", x"0c74", x"0c74", x"0c74", x"0c75", x"0c75", x"0c75", x"0c75", x"0c75", x"0c75", x"0c76", x"0c76", x"0c76", x"0c76", x"0c76", x"0c76", x"0c77", x"0c77", x"0c77", x"0c77", x"0c77", x"0c78", x"0c78", x"0c78", x"0c78", x"0c78", x"0c78", x"0c79", x"0c79", x"0c79", x"0c79", x"0c79", x"0c79", x"0c7a", x"0c7a", x"0c7a", x"0c7a", x"0c7a", x"0c7a", x"0c7b", x"0c7b", x"0c7b", x"0c7b", x"0c7b", x"0c7b", x"0c7c", x"0c7c", x"0c7c", x"0c7c", x"0c7c", x"0c7c", x"0c7d", x"0c7d", x"0c7d", x"0c7d", x"0c7d", x"0c7e", x"0c7e", x"0c7e", x"0c7e", x"0c7e", x"0c7e", x"0c7f", x"0c7f", x"0c7f", x"0c7f", x"0c7f", x"0c7f", x"0c80", x"0c80", x"0c80", x"0c80", x"0c80", x"0c80", x"0c81", x"0c81", x"0c81", x"0c81", x"0c81", x"0c81", x"0c82", x"0c82", x"0c82", x"0c82", x"0c82", x"0c82", x"0c83", x"0c83", x"0c83", x"0c83", x"0c83", x"0c83", x"0c84", x"0c84", x"0c84", x"0c84", x"0c84", x"0c85", x"0c85", x"0c85", x"0c85", x"0c85", x"0c85", x"0c86", x"0c86", x"0c86", x"0c86", x"0c86", x"0c86", x"0c87", x"0c87", x"0c87", x"0c87", x"0c87", x"0c87", x"0c88", x"0c88", x"0c88", x"0c88", x"0c88", x"0c88", x"0c89", x"0c89", x"0c89", x"0c89", x"0c89", x"0c89", x"0c8a", x"0c8a", x"0c8a", x"0c8a", x"0c8a", x"0c8a", x"0c8b", x"0c8b", x"0c8b", x"0c8b", x"0c8b", x"0c8b", x"0c8c", x"0c8c", x"0c8c", x"0c8c", x"0c8c", x"0c8c", x"0c8d", x"0c8d", x"0c8d", x"0c8d", x"0c8d", x"0c8d", x"0c8e", x"0c8e", x"0c8e", x"0c8e", x"0c8e", x"0c8e", x"0c8f", x"0c8f", x"0c8f", x"0c8f", x"0c8f", x"0c90", x"0c90", x"0c90", x"0c90", x"0c90", x"0c90", x"0c91", x"0c91", x"0c91", x"0c91", x"0c91", x"0c91", x"0c92", x"0c92", x"0c92", x"0c92", x"0c92", x"0c92", x"0c93", x"0c93", x"0c93", x"0c93", x"0c93", x"0c93", x"0c94", x"0c94", x"0c94", x"0c94", x"0c94", x"0c94", x"0c95", x"0c95", x"0c95", x"0c95", x"0c95", x"0c95", x"0c96", x"0c96", x"0c96", x"0c96", x"0c96", x"0c96", x"0c97", x"0c97", x"0c97", x"0c97", x"0c97", x"0c97", x"0c98", x"0c98", x"0c98", x"0c98", x"0c98", x"0c98", x"0c99", x"0c99", x"0c99", x"0c99", x"0c99", x"0c99", x"0c9a", x"0c9a", x"0c9a", x"0c9a", x"0c9a", x"0c9a", x"0c9b", x"0c9b", x"0c9b", x"0c9b", x"0c9b", x"0c9b", x"0c9c", x"0c9c", x"0c9c", x"0c9c", x"0c9c", x"0c9c", x"0c9d", x"0c9d", x"0c9d", x"0c9d", x"0c9d", x"0c9d", x"0c9e", x"0c9e", x"0c9e", x"0c9e", x"0c9e", x"0c9e", x"0c9f", x"0c9f", x"0c9f", x"0c9f", x"0c9f", x"0c9f", x"0ca0", x"0ca0", x"0ca0", x"0ca0", x"0ca0", x"0ca0", x"0ca1", x"0ca1", x"0ca1", x"0ca1", x"0ca1", x"0ca1", x"0ca2", x"0ca2", x"0ca2", x"0ca2", x"0ca2", x"0ca2", x"0ca3", x"0ca3", x"0ca3", x"0ca3", x"0ca3", x"0ca3", x"0ca4", x"0ca4", x"0ca4", x"0ca4", x"0ca4", x"0ca4", x"0ca5", x"0ca5", x"0ca5", x"0ca5", x"0ca5", x"0ca5", x"0ca6", x"0ca6", x"0ca6", x"0ca6", x"0ca6", x"0ca6", x"0ca7", x"0ca7", x"0ca7", x"0ca7", x"0ca7", x"0ca7", x"0ca8", x"0ca8", x"0ca8", x"0ca8", x"0ca8", x"0ca8", x"0ca9", x"0ca9", x"0ca9", x"0ca9", x"0ca9", x"0ca9", x"0caa", x"0caa", x"0caa", x"0caa", x"0caa", x"0caa", x"0cab", x"0cab", x"0cab", x"0cab", x"0cab", x"0cab", x"0cab", x"0cac", x"0cac", x"0cac", x"0cac", x"0cac", x"0cac", x"0cad", x"0cad", x"0cad", x"0cad", x"0cad", x"0cad", x"0cae", x"0cae", x"0cae", x"0cae", x"0cae", x"0cae", x"0caf", x"0caf", x"0caf", x"0caf", x"0caf", x"0caf", x"0cb0", x"0cb0", x"0cb0", x"0cb0", x"0cb0", x"0cb0", x"0cb1", x"0cb1", x"0cb1", x"0cb1", x"0cb1", x"0cb1", x"0cb2", x"0cb2", x"0cb2", x"0cb2", x"0cb2", x"0cb2", x"0cb3", x"0cb3", x"0cb3", x"0cb3", x"0cb3", x"0cb3", x"0cb4", x"0cb4", x"0cb4", x"0cb4", x"0cb4", x"0cb4", x"0cb5", x"0cb5", x"0cb5", x"0cb5", x"0cb5", x"0cb5", x"0cb5", x"0cb6", x"0cb6", x"0cb6", x"0cb6", x"0cb6", x"0cb6", x"0cb7", x"0cb7", x"0cb7", x"0cb7", x"0cb7", x"0cb7", x"0cb8", x"0cb8", x"0cb8", x"0cb8", x"0cb8", x"0cb8", x"0cb9", x"0cb9", x"0cb9", x"0cb9", x"0cb9", x"0cb9", x"0cba", x"0cba", x"0cba", x"0cba", x"0cba", x"0cba", x"0cbb", x"0cbb", x"0cbb", x"0cbb", x"0cbb", x"0cbb", x"0cbc", x"0cbc", x"0cbc", x"0cbc", x"0cbc", x"0cbc", x"0cbc", x"0cbd", x"0cbd", x"0cbd", x"0cbd", x"0cbd", x"0cbd", x"0cbe", x"0cbe", x"0cbe", x"0cbe", x"0cbe", x"0cbe", x"0cbf", x"0cbf", x"0cbf", x"0cbf", x"0cbf", x"0cbf", x"0cc0", x"0cc0", x"0cc0", x"0cc0", x"0cc0", x"0cc0", x"0cc1", x"0cc1", x"0cc1", x"0cc1", x"0cc1", x"0cc1", x"0cc1", x"0cc2", x"0cc2", x"0cc2", x"0cc2", x"0cc2", x"0cc2", x"0cc3", x"0cc3", x"0cc3", x"0cc3", x"0cc3", x"0cc3", x"0cc4", x"0cc4", x"0cc4", x"0cc4", x"0cc4", x"0cc4", x"0cc5", x"0cc5", x"0cc5", x"0cc5", x"0cc5", x"0cc5", x"0cc6", x"0cc6", x"0cc6", x"0cc6", x"0cc6", x"0cc6", x"0cc6", x"0cc7", x"0cc7", x"0cc7", x"0cc7", x"0cc7", x"0cc7", x"0cc8", x"0cc8", x"0cc8", x"0cc8", x"0cc8", x"0cc8", x"0cc9", x"0cc9", x"0cc9", x"0cc9", x"0cc9", x"0cc9", x"0cca", x"0cca", x"0cca", x"0cca", x"0cca", x"0cca", x"0cca", x"0ccb", x"0ccb", x"0ccb", x"0ccb", x"0ccb", x"0ccb", x"0ccc", x"0ccc", x"0ccc", x"0ccc", x"0ccc", x"0ccc", x"0ccd", x"0ccd", x"0ccd", x"0ccd", x"0ccd", x"0ccd", x"0cce", x"0cce", x"0cce", x"0cce", x"0cce", x"0cce", x"0cce", x"0ccf", x"0ccf", x"0ccf", x"0ccf", x"0ccf", x"0ccf", x"0cd0", x"0cd0", x"0cd0", x"0cd0", x"0cd0", x"0cd0", x"0cd1", x"0cd1", x"0cd1", x"0cd1", x"0cd1", x"0cd1", x"0cd2", x"0cd2", x"0cd2", x"0cd2", x"0cd2", x"0cd2", x"0cd2", x"0cd3", x"0cd3", x"0cd3", x"0cd3", x"0cd3", x"0cd3", x"0cd4", x"0cd4", x"0cd4", x"0cd4", x"0cd4", x"0cd4", x"0cd5", x"0cd5", x"0cd5", x"0cd5", x"0cd5", x"0cd5", x"0cd5", x"0cd6", x"0cd6", x"0cd6", x"0cd6", x"0cd6", x"0cd6", x"0cd7", x"0cd7", x"0cd7", x"0cd7", x"0cd7", x"0cd7", x"0cd8", x"0cd8", x"0cd8", x"0cd8", x"0cd8", x"0cd8", x"0cd8", x"0cd9", x"0cd9", x"0cd9", x"0cd9", x"0cd9", x"0cd9", x"0cda", x"0cda", x"0cda", x"0cda", x"0cda", x"0cda", x"0cdb", x"0cdb", x"0cdb", x"0cdb", x"0cdb", x"0cdb", x"0cdb", x"0cdc", x"0cdc", x"0cdc", x"0cdc", x"0cdc", x"0cdc", x"0cdd", x"0cdd", x"0cdd", x"0cdd", x"0cdd", x"0cdd", x"0cde", x"0cde", x"0cde", x"0cde", x"0cde", x"0cde", x"0cde", x"0cdf", x"0cdf", x"0cdf", x"0cdf", x"0cdf", x"0cdf", x"0ce0", x"0ce0", x"0ce0", x"0ce0", x"0ce0", x"0ce0", x"0ce1", x"0ce1", x"0ce1", x"0ce1", x"0ce1", x"0ce1", x"0ce1", x"0ce2", x"0ce2", x"0ce2", x"0ce2", x"0ce2", x"0ce2", x"0ce3", x"0ce3", x"0ce3", x"0ce3", x"0ce3", x"0ce3", x"0ce4", x"0ce4", x"0ce4", x"0ce4", x"0ce4", x"0ce4", x"0ce4", x"0ce5", x"0ce5", x"0ce5", x"0ce5", x"0ce5", x"0ce5", x"0ce6", x"0ce6", x"0ce6", x"0ce6", x"0ce6", x"0ce6", x"0ce6", x"0ce7", x"0ce7", x"0ce7", x"0ce7", x"0ce7", x"0ce7", x"0ce8", x"0ce8", x"0ce8", x"0ce8", x"0ce8", x"0ce8", x"0ce8", x"0ce9", x"0ce9", x"0ce9", x"0ce9", x"0ce9", x"0ce9", x"0cea", x"0cea", x"0cea", x"0cea", x"0cea", x"0cea", x"0ceb", x"0ceb", x"0ceb", x"0ceb", x"0ceb", x"0ceb", x"0ceb", x"0cec", x"0cec", x"0cec", x"0cec", x"0cec", x"0cec", x"0ced", x"0ced", x"0ced", x"0ced", x"0ced", x"0ced", x"0ced", x"0cee", x"0cee", x"0cee", x"0cee", x"0cee", x"0cee", x"0cef", x"0cef", x"0cef", x"0cef", x"0cef", x"0cef", x"0cef", x"0cf0", x"0cf0", x"0cf0", x"0cf0", x"0cf0", x"0cf0", x"0cf1", x"0cf1", x"0cf1", x"0cf1", x"0cf1", x"0cf1", x"0cf1", x"0cf2", x"0cf2", x"0cf2", x"0cf2", x"0cf2", x"0cf2", x"0cf3", x"0cf3", x"0cf3", x"0cf3", x"0cf3", x"0cf3", x"0cf3", x"0cf4", x"0cf4", x"0cf4", x"0cf4", x"0cf4", x"0cf4", x"0cf5", x"0cf5", x"0cf5", x"0cf5", x"0cf5", x"0cf5", x"0cf5", x"0cf6", x"0cf6", x"0cf6", x"0cf6", x"0cf6", x"0cf6", x"0cf7", x"0cf7", x"0cf7", x"0cf7", x"0cf7", x"0cf7", x"0cf7", x"0cf8", x"0cf8", x"0cf8", x"0cf8", x"0cf8", x"0cf8", x"0cf9", x"0cf9", x"0cf9", x"0cf9", x"0cf9", x"0cf9", x"0cf9", x"0cfa", x"0cfa", x"0cfa", x"0cfa", x"0cfa", x"0cfa", x"0cfb", x"0cfb", x"0cfb", x"0cfb", x"0cfb", x"0cfb", x"0cfb", x"0cfc", x"0cfc", x"0cfc", x"0cfc", x"0cfc", x"0cfc", x"0cfd", x"0cfd", x"0cfd", x"0cfd", x"0cfd", x"0cfd", x"0cfd", x"0cfe", x"0cfe", x"0cfe", x"0cfe", x"0cfe", x"0cfe", x"0cff", x"0cff", x"0cff", x"0cff", x"0cff", x"0cff", x"0cff", x"0d00", x"0d00", x"0d00", x"0d00", x"0d00", x"0d00", x"0d00", x"0d01", x"0d01", x"0d01", x"0d01", x"0d01", x"0d01", x"0d02", x"0d02", x"0d02", x"0d02", x"0d02", x"0d02", x"0d02", x"0d03", x"0d03", x"0d03", x"0d03", x"0d03", x"0d03", x"0d04", x"0d04", x"0d04", x"0d04", x"0d04", x"0d04", x"0d04", x"0d05", x"0d05", x"0d05", x"0d05", x"0d05", x"0d05", x"0d06", x"0d06", x"0d06", x"0d06", x"0d06", x"0d06", x"0d06", x"0d07", x"0d07", x"0d07", x"0d07", x"0d07", x"0d07", x"0d07", x"0d08", x"0d08", x"0d08", x"0d08", x"0d08", x"0d08", x"0d09", x"0d09", x"0d09", x"0d09", x"0d09", x"0d09", x"0d09", x"0d0a", x"0d0a", x"0d0a", x"0d0a", x"0d0a", x"0d0a", x"0d0a", x"0d0b", x"0d0b", x"0d0b", x"0d0b", x"0d0b", x"0d0b", x"0d0c", x"0d0c", x"0d0c", x"0d0c", x"0d0c", x"0d0c", x"0d0c", x"0d0d", x"0d0d", x"0d0d", x"0d0d", x"0d0d", x"0d0d", x"0d0d", x"0d0e", x"0d0e", x"0d0e", x"0d0e", x"0d0e", x"0d0e", x"0d0f", x"0d0f", x"0d0f", x"0d0f", x"0d0f", x"0d0f", x"0d0f", x"0d10", x"0d10", x"0d10", x"0d10", x"0d10", x"0d10", x"0d10", x"0d11", x"0d11", x"0d11", x"0d11", x"0d11", x"0d11", x"0d12", x"0d12", x"0d12", x"0d12", x"0d12", x"0d12", x"0d12", x"0d13", x"0d13", x"0d13", x"0d13", x"0d13", x"0d13", x"0d13", x"0d14", x"0d14", x"0d14", x"0d14", x"0d14", x"0d14", x"0d15", x"0d15", x"0d15", x"0d15", x"0d15", x"0d15", x"0d15", x"0d16", x"0d16", x"0d16", x"0d16", x"0d16", x"0d16", x"0d16", x"0d17", x"0d17", x"0d17", x"0d17", x"0d17", x"0d17", x"0d17", x"0d18", x"0d18", x"0d18", x"0d18", x"0d18", x"0d18", x"0d19", x"0d19", x"0d19", x"0d19", x"0d19", x"0d19", x"0d19", x"0d1a", x"0d1a", x"0d1a", x"0d1a", x"0d1a", x"0d1a", x"0d1a", x"0d1b", x"0d1b", x"0d1b", x"0d1b", x"0d1b", x"0d1b", x"0d1b", x"0d1c", x"0d1c", x"0d1c", x"0d1c", x"0d1c", x"0d1c", x"0d1d", x"0d1d", x"0d1d", x"0d1d", x"0d1d", x"0d1d", x"0d1d", x"0d1e", x"0d1e", x"0d1e", x"0d1e", x"0d1e", x"0d1e", x"0d1e", x"0d1f", x"0d1f", x"0d1f", x"0d1f", x"0d1f", x"0d1f", x"0d1f", x"0d20", x"0d20", x"0d20", x"0d20", x"0d20", x"0d20", x"0d20", x"0d21", x"0d21", x"0d21", x"0d21", x"0d21", x"0d21", x"0d22", x"0d22", x"0d22", x"0d22", x"0d22", x"0d22", x"0d22", x"0d23", x"0d23", x"0d23", x"0d23", x"0d23", x"0d23", x"0d23", x"0d24", x"0d24", x"0d24", x"0d24", x"0d24", x"0d24", x"0d24", x"0d25", x"0d25", x"0d25", x"0d25", x"0d25", x"0d25", x"0d25", x"0d26", x"0d26", x"0d26", x"0d26", x"0d26", x"0d26", x"0d27", x"0d27", x"0d27", x"0d27", x"0d27", x"0d27", x"0d27", x"0d28", x"0d28", x"0d28", x"0d28", x"0d28", x"0d28", x"0d28", x"0d29", x"0d29", x"0d29", x"0d29", x"0d29", x"0d29", x"0d29", x"0d2a", x"0d2a", x"0d2a", x"0d2a", x"0d2a", x"0d2a", x"0d2a", x"0d2b", x"0d2b", x"0d2b", x"0d2b", x"0d2b", x"0d2b", x"0d2b", x"0d2c", x"0d2c", x"0d2c", x"0d2c", x"0d2c", x"0d2c", x"0d2c", x"0d2d", x"0d2d", x"0d2d", x"0d2d", x"0d2d", x"0d2d", x"0d2d", x"0d2e", x"0d2e", x"0d2e", x"0d2e", x"0d2e", x"0d2e", x"0d2f", x"0d2f", x"0d2f", x"0d2f", x"0d2f", x"0d2f", x"0d2f", x"0d30", x"0d30", x"0d30", x"0d30", x"0d30", x"0d30", x"0d30", x"0d31", x"0d31", x"0d31", x"0d31", x"0d31", x"0d31", x"0d31", x"0d32", x"0d32", x"0d32", x"0d32", x"0d32", x"0d32", x"0d32", x"0d33", x"0d33", x"0d33", x"0d33", x"0d33", x"0d33", x"0d33", x"0d34", x"0d34", x"0d34", x"0d34", x"0d34", x"0d34", x"0d34", x"0d35", x"0d35", x"0d35", x"0d35", x"0d35", x"0d35", x"0d35", x"0d36", x"0d36", x"0d36", x"0d36", x"0d36", x"0d36", x"0d36", x"0d37", x"0d37", x"0d37", x"0d37", x"0d37", x"0d37", x"0d37", x"0d38", x"0d38", x"0d38", x"0d38", x"0d38", x"0d38", x"0d38", x"0d39", x"0d39", x"0d39", x"0d39", x"0d39", x"0d39", x"0d39", x"0d3a", x"0d3a", x"0d3a", x"0d3a", x"0d3a", x"0d3a", x"0d3a", x"0d3b", x"0d3b", x"0d3b", x"0d3b", x"0d3b", x"0d3b", x"0d3b", x"0d3c", x"0d3c", x"0d3c", x"0d3c", x"0d3c", x"0d3c", x"0d3c", x"0d3d", x"0d3d", x"0d3d", x"0d3d", x"0d3d", x"0d3d", x"0d3d", x"0d3e", x"0d3e", x"0d3e", x"0d3e", x"0d3e", x"0d3e", x"0d3e", x"0d3f", x"0d3f", x"0d3f", x"0d3f", x"0d3f", x"0d3f", x"0d3f", x"0d40", x"0d40", x"0d40", x"0d40", x"0d40", x"0d40", x"0d40", x"0d41", x"0d41", x"0d41", x"0d41", x"0d41", x"0d41", x"0d41", x"0d42", x"0d42", x"0d42", x"0d42", x"0d42", x"0d42", x"0d42", x"0d43", x"0d43", x"0d43", x"0d43", x"0d43", x"0d43", x"0d43", x"0d44", x"0d44", x"0d44", x"0d44", x"0d44", x"0d44", x"0d44", x"0d45", x"0d45", x"0d45", x"0d45", x"0d45", x"0d45", x"0d45", x"0d46", x"0d46", x"0d46", x"0d46", x"0d46", x"0d46", x"0d46", x"0d47", x"0d47", x"0d47", x"0d47", x"0d47", x"0d47", x"0d47", x"0d48", x"0d48", x"0d48", x"0d48", x"0d48", x"0d48", x"0d48", x"0d49", x"0d49", x"0d49", x"0d49", x"0d49", x"0d49", x"0d49", x"0d49", x"0d4a", x"0d4a", x"0d4a", x"0d4a", x"0d4a", x"0d4a", x"0d4a", x"0d4b", x"0d4b", x"0d4b", x"0d4b", x"0d4b", x"0d4b", x"0d4b", x"0d4c", x"0d4c", x"0d4c", x"0d4c", x"0d4c", x"0d4c", x"0d4c", x"0d4d", x"0d4d", x"0d4d", x"0d4d", x"0d4d", x"0d4d", x"0d4d", x"0d4e", x"0d4e", x"0d4e", x"0d4e", x"0d4e", x"0d4e", x"0d4e", x"0d4f", x"0d4f", x"0d4f", x"0d4f", x"0d4f", x"0d4f", x"0d4f", x"0d50", x"0d50", x"0d50", x"0d50", x"0d50", x"0d50", x"0d50", x"0d50", x"0d51", x"0d51", x"0d51", x"0d51", x"0d51", x"0d51", x"0d51", x"0d52", x"0d52", x"0d52", x"0d52", x"0d52", x"0d52", x"0d52", x"0d53", x"0d53", x"0d53", x"0d53", x"0d53", x"0d53", x"0d53", x"0d54", x"0d54", x"0d54", x"0d54", x"0d54", x"0d54", x"0d54", x"0d55", x"0d55", x"0d55", x"0d55", x"0d55", x"0d55", x"0d55", x"0d55", x"0d56", x"0d56", x"0d56", x"0d56", x"0d56", x"0d56", x"0d56", x"0d57", x"0d57", x"0d57", x"0d57", x"0d57", x"0d57", x"0d57", x"0d58", x"0d58", x"0d58", x"0d58", x"0d58", x"0d58", x"0d58", x"0d59", x"0d59", x"0d59", x"0d59", x"0d59", x"0d59", x"0d59", x"0d5a", x"0d5a", x"0d5a", x"0d5a", x"0d5a", x"0d5a", x"0d5a", x"0d5a", x"0d5b", x"0d5b", x"0d5b", x"0d5b", x"0d5b", x"0d5b", x"0d5b", x"0d5c", x"0d5c", x"0d5c", x"0d5c", x"0d5c", x"0d5c", x"0d5c", x"0d5d", x"0d5d", x"0d5d", x"0d5d", x"0d5d", x"0d5d", x"0d5d", x"0d5d", x"0d5e", x"0d5e", x"0d5e", x"0d5e", x"0d5e", x"0d5e", x"0d5e", x"0d5f", x"0d5f", x"0d5f", x"0d5f", x"0d5f", x"0d5f", x"0d5f", x"0d60", x"0d60", x"0d60", x"0d60", x"0d60", x"0d60", x"0d60", x"0d61", x"0d61", x"0d61", x"0d61", x"0d61", x"0d61", x"0d61", x"0d61", x"0d62", x"0d62", x"0d62", x"0d62", x"0d62", x"0d62", x"0d62", x"0d63", x"0d63", x"0d63", x"0d63", x"0d63", x"0d63", x"0d63", x"0d64", x"0d64", x"0d64", x"0d64", x"0d64", x"0d64", x"0d64", x"0d64", x"0d65", x"0d65", x"0d65", x"0d65", x"0d65", x"0d65", x"0d65", x"0d66", x"0d66", x"0d66", x"0d66", x"0d66", x"0d66", x"0d66", x"0d67", x"0d67", x"0d67", x"0d67", x"0d67", x"0d67", x"0d67", x"0d67", x"0d68", x"0d68", x"0d68", x"0d68", x"0d68", x"0d68", x"0d68", x"0d69", x"0d69", x"0d69", x"0d69", x"0d69", x"0d69", x"0d69", x"0d69", x"0d6a", x"0d6a", x"0d6a", x"0d6a", x"0d6a", x"0d6a", x"0d6a", x"0d6b", x"0d6b", x"0d6b", x"0d6b", x"0d6b", x"0d6b", x"0d6b", x"0d6c", x"0d6c", x"0d6c", x"0d6c", x"0d6c", x"0d6c", x"0d6c", x"0d6c", x"0d6d", x"0d6d", x"0d6d", x"0d6d", x"0d6d", x"0d6d", x"0d6d", x"0d6e", x"0d6e", x"0d6e", x"0d6e", x"0d6e", x"0d6e", x"0d6e", x"0d6e", x"0d6f", x"0d6f", x"0d6f", x"0d6f", x"0d6f", x"0d6f", x"0d6f", x"0d70", x"0d70", x"0d70", x"0d70", x"0d70", x"0d70", x"0d70", x"0d70", x"0d71", x"0d71", x"0d71", x"0d71", x"0d71", x"0d71", x"0d71", x"0d72", x"0d72", x"0d72", x"0d72", x"0d72", x"0d72", x"0d72", x"0d73", x"0d73", x"0d73", x"0d73", x"0d73", x"0d73", x"0d73", x"0d73", x"0d74", x"0d74", x"0d74", x"0d74", x"0d74", x"0d74", x"0d74", x"0d75", x"0d75", x"0d75", x"0d75", x"0d75", x"0d75", x"0d75", x"0d75", x"0d76", x"0d76", x"0d76", x"0d76", x"0d76", x"0d76", x"0d76", x"0d77", x"0d77", x"0d77", x"0d77", x"0d77", x"0d77", x"0d77", x"0d77", x"0d78", x"0d78", x"0d78", x"0d78", x"0d78", x"0d78", x"0d78", x"0d79", x"0d79", x"0d79", x"0d79", x"0d79", x"0d79", x"0d79", x"0d79", x"0d7a", x"0d7a", x"0d7a", x"0d7a", x"0d7a", x"0d7a", x"0d7a", x"0d7a", x"0d7b", x"0d7b", x"0d7b", x"0d7b", x"0d7b", x"0d7b", x"0d7b", x"0d7c", x"0d7c", x"0d7c", x"0d7c", x"0d7c", x"0d7c", x"0d7c", x"0d7c", x"0d7d", x"0d7d", x"0d7d", x"0d7d", x"0d7d", x"0d7d", x"0d7d", x"0d7e", x"0d7e", x"0d7e", x"0d7e", x"0d7e", x"0d7e", x"0d7e", x"0d7e", x"0d7f", x"0d7f", x"0d7f", x"0d7f", x"0d7f", x"0d7f", x"0d7f", x"0d80", x"0d80", x"0d80", x"0d80", x"0d80", x"0d80", x"0d80", x"0d80", x"0d81", x"0d81", x"0d81", x"0d81", x"0d81", x"0d81", x"0d81", x"0d81", x"0d82", x"0d82", x"0d82", x"0d82", x"0d82", x"0d82", x"0d82", x"0d83", x"0d83", x"0d83", x"0d83", x"0d83", x"0d83", x"0d83", x"0d83", x"0d84", x"0d84", x"0d84", x"0d84", x"0d84", x"0d84", x"0d84", x"0d85", x"0d85", x"0d85", x"0d85", x"0d85", x"0d85", x"0d85", x"0d85", x"0d86", x"0d86", x"0d86", x"0d86", x"0d86", x"0d86", x"0d86", x"0d86", x"0d87", x"0d87", x"0d87", x"0d87", x"0d87", x"0d87", x"0d87", x"0d88", x"0d88", x"0d88", x"0d88", x"0d88", x"0d88", x"0d88", x"0d88", x"0d89", x"0d89", x"0d89", x"0d89", x"0d89", x"0d89", x"0d89", x"0d89", x"0d8a", x"0d8a", x"0d8a", x"0d8a", x"0d8a", x"0d8a", x"0d8a", x"0d8a", x"0d8b", x"0d8b", x"0d8b", x"0d8b", x"0d8b", x"0d8b", x"0d8b", x"0d8c", x"0d8c", x"0d8c", x"0d8c", x"0d8c", x"0d8c", x"0d8c", x"0d8c", x"0d8d", x"0d8d", x"0d8d", x"0d8d", x"0d8d", x"0d8d", x"0d8d", x"0d8d", x"0d8e", x"0d8e", x"0d8e", x"0d8e", x"0d8e", x"0d8e", x"0d8e", x"0d8f", x"0d8f", x"0d8f", x"0d8f", x"0d8f", x"0d8f", x"0d8f", x"0d8f", x"0d90", x"0d90", x"0d90", x"0d90", x"0d90", x"0d90", x"0d90", x"0d90", x"0d91", x"0d91", x"0d91", x"0d91", x"0d91", x"0d91", x"0d91", x"0d91", x"0d92", x"0d92", x"0d92", x"0d92", x"0d92", x"0d92", x"0d92", x"0d93", x"0d93", x"0d93", x"0d93", x"0d93", x"0d93", x"0d93", x"0d93", x"0d94", x"0d94", x"0d94", x"0d94", x"0d94", x"0d94", x"0d94", x"0d94", x"0d95", x"0d95", x"0d95", x"0d95", x"0d95", x"0d95", x"0d95", x"0d95", x"0d96", x"0d96", x"0d96", x"0d96", x"0d96", x"0d96", x"0d96", x"0d96", x"0d97", x"0d97", x"0d97", x"0d97", x"0d97", x"0d97", x"0d97", x"0d97", x"0d98", x"0d98", x"0d98", x"0d98", x"0d98", x"0d98", x"0d98", x"0d99", x"0d99", x"0d99", x"0d99", x"0d99", x"0d99", x"0d99", x"0d99", x"0d9a", x"0d9a", x"0d9a", x"0d9a", x"0d9a", x"0d9a", x"0d9a", x"0d9a", x"0d9b", x"0d9b", x"0d9b", x"0d9b", x"0d9b", x"0d9b", x"0d9b", x"0d9b", x"0d9c", x"0d9c", x"0d9c", x"0d9c", x"0d9c", x"0d9c", x"0d9c", x"0d9c", x"0d9d", x"0d9d", x"0d9d", x"0d9d", x"0d9d", x"0d9d", x"0d9d", x"0d9d", x"0d9e", x"0d9e", x"0d9e", x"0d9e", x"0d9e", x"0d9e", x"0d9e", x"0d9e", x"0d9f", x"0d9f", x"0d9f", x"0d9f", x"0d9f", x"0d9f", x"0d9f", x"0d9f", x"0da0", x"0da0", x"0da0", x"0da0", x"0da0", x"0da0", x"0da0", x"0da0", x"0da1", x"0da1", x"0da1", x"0da1", x"0da1", x"0da1", x"0da1", x"0da2", x"0da2", x"0da2", x"0da2", x"0da2", x"0da2", x"0da2", x"0da2", x"0da3", x"0da3", x"0da3", x"0da3", x"0da3", x"0da3", x"0da3", x"0da3", x"0da4", x"0da4", x"0da4", x"0da4", x"0da4", x"0da4", x"0da4", x"0da4", x"0da5", x"0da5", x"0da5", x"0da5", x"0da5", x"0da5", x"0da5", x"0da5", x"0da6", x"0da6", x"0da6", x"0da6", x"0da6", x"0da6", x"0da6", x"0da6", x"0da7", x"0da7", x"0da7", x"0da7", x"0da7", x"0da7", x"0da7", x"0da7", x"0da8", x"0da8", x"0da8", x"0da8", x"0da8", x"0da8", x"0da8", x"0da8", x"0da9", x"0da9", x"0da9", x"0da9", x"0da9", x"0da9", x"0da9", x"0da9", x"0daa", x"0daa", x"0daa", x"0daa", x"0daa", x"0daa", x"0daa", x"0daa", x"0dab", x"0dab", x"0dab", x"0dab", x"0dab", x"0dab", x"0dab", x"0dab", x"0dac", x"0dac", x"0dac", x"0dac", x"0dac", x"0dac", x"0dac", x"0dac", x"0dad", x"0dad", x"0dad", x"0dad", x"0dad", x"0dad", x"0dad", x"0dad", x"0dad", x"0dae", x"0dae", x"0dae", x"0dae", x"0dae", x"0dae", x"0dae", x"0dae", x"0daf", x"0daf", x"0daf", x"0daf", x"0daf", x"0daf", x"0daf", x"0daf", x"0db0", x"0db0", x"0db0", x"0db0", x"0db0", x"0db0", x"0db0", x"0db0", x"0db1", x"0db1", x"0db1", x"0db1", x"0db1", x"0db1", x"0db1", x"0db1", x"0db2", x"0db2", x"0db2", x"0db2", x"0db2", x"0db2", x"0db2", x"0db2", x"0db3", x"0db3", x"0db3", x"0db3", x"0db3", x"0db3", x"0db3", x"0db3", x"0db4", x"0db4", x"0db4", x"0db4", x"0db4", x"0db4", x"0db4", x"0db4", x"0db5", x"0db5", x"0db5", x"0db5", x"0db5", x"0db5", x"0db5", x"0db5", x"0db5", x"0db6", x"0db6", x"0db6", x"0db6", x"0db6", x"0db6", x"0db6", x"0db6", x"0db7", x"0db7", x"0db7", x"0db7", x"0db7", x"0db7", x"0db7", x"0db7", x"0db8", x"0db8", x"0db8", x"0db8", x"0db8", x"0db8", x"0db8", x"0db8", x"0db9", x"0db9", x"0db9", x"0db9", x"0db9", x"0db9", x"0db9", x"0db9", x"0dba", x"0dba", x"0dba", x"0dba", x"0dba", x"0dba", x"0dba", x"0dba", x"0dba", x"0dbb", x"0dbb", x"0dbb", x"0dbb", x"0dbb", x"0dbb", x"0dbb", x"0dbb", x"0dbc", x"0dbc", x"0dbc", x"0dbc", x"0dbc", x"0dbc", x"0dbc", x"0dbc", x"0dbd", x"0dbd", x"0dbd", x"0dbd", x"0dbd", x"0dbd", x"0dbd", x"0dbd", x"0dbe", x"0dbe", x"0dbe", x"0dbe", x"0dbe", x"0dbe", x"0dbe", x"0dbe", x"0dbe", x"0dbf", x"0dbf", x"0dbf", x"0dbf", x"0dbf", x"0dbf", x"0dbf", x"0dbf", x"0dc0", x"0dc0", x"0dc0", x"0dc0", x"0dc0", x"0dc0", x"0dc0", x"0dc0", x"0dc1", x"0dc1", x"0dc1", x"0dc1", x"0dc1", x"0dc1", x"0dc1", x"0dc1", x"0dc2", x"0dc2", x"0dc2", x"0dc2", x"0dc2", x"0dc2", x"0dc2", x"0dc2", x"0dc2", x"0dc3", x"0dc3", x"0dc3", x"0dc3", x"0dc3", x"0dc3", x"0dc3", x"0dc3", x"0dc4", x"0dc4", x"0dc4", x"0dc4", x"0dc4", x"0dc4", x"0dc4", x"0dc4", x"0dc5", x"0dc5", x"0dc5", x"0dc5", x"0dc5", x"0dc5", x"0dc5", x"0dc5", x"0dc5", x"0dc6", x"0dc6", x"0dc6", x"0dc6", x"0dc6", x"0dc6", x"0dc6", x"0dc6", x"0dc7", x"0dc7", x"0dc7", x"0dc7", x"0dc7", x"0dc7", x"0dc7", x"0dc7", x"0dc7", x"0dc8", x"0dc8", x"0dc8", x"0dc8", x"0dc8", x"0dc8", x"0dc8", x"0dc8", x"0dc9", x"0dc9", x"0dc9", x"0dc9", x"0dc9", x"0dc9", x"0dc9", x"0dc9", x"0dca", x"0dca", x"0dca", x"0dca", x"0dca", x"0dca", x"0dca", x"0dca", x"0dca", x"0dcb", x"0dcb", x"0dcb", x"0dcb", x"0dcb", x"0dcb", x"0dcb", x"0dcb", x"0dcc", x"0dcc", x"0dcc", x"0dcc", x"0dcc", x"0dcc", x"0dcc", x"0dcc", x"0dcc", x"0dcd", x"0dcd", x"0dcd", x"0dcd", x"0dcd", x"0dcd", x"0dcd", x"0dcd", x"0dce", x"0dce", x"0dce", x"0dce", x"0dce", x"0dce", x"0dce", x"0dce", x"0dce", x"0dcf", x"0dcf", x"0dcf", x"0dcf", x"0dcf", x"0dcf", x"0dcf", x"0dcf", x"0dd0", x"0dd0", x"0dd0", x"0dd0", x"0dd0", x"0dd0", x"0dd0", x"0dd0", x"0dd1", x"0dd1", x"0dd1", x"0dd1", x"0dd1", x"0dd1", x"0dd1", x"0dd1", x"0dd1", x"0dd2", x"0dd2", x"0dd2", x"0dd2", x"0dd2", x"0dd2", x"0dd2", x"0dd2", x"0dd2", x"0dd3", x"0dd3", x"0dd3", x"0dd3", x"0dd3", x"0dd3", x"0dd3", x"0dd3", x"0dd4", x"0dd4", x"0dd4", x"0dd4", x"0dd4", x"0dd4", x"0dd4", x"0dd4", x"0dd4", x"0dd5", x"0dd5", x"0dd5", x"0dd5", x"0dd5", x"0dd5", x"0dd5", x"0dd5", x"0dd6", x"0dd6", x"0dd6", x"0dd6", x"0dd6", x"0dd6", x"0dd6", x"0dd6", x"0dd6", x"0dd7", x"0dd7", x"0dd7", x"0dd7", x"0dd7", x"0dd7", x"0dd7", x"0dd7", x"0dd8", x"0dd8", x"0dd8", x"0dd8", x"0dd8", x"0dd8", x"0dd8", x"0dd8", x"0dd8", x"0dd9", x"0dd9", x"0dd9", x"0dd9", x"0dd9", x"0dd9", x"0dd9", x"0dd9", x"0dda", x"0dda", x"0dda", x"0dda", x"0dda", x"0dda", x"0dda", x"0dda", x"0dda", x"0ddb", x"0ddb", x"0ddb", x"0ddb", x"0ddb", x"0ddb", x"0ddb", x"0ddb", x"0ddb", x"0ddc", x"0ddc", x"0ddc", x"0ddc", x"0ddc", x"0ddc", x"0ddc", x"0ddc", x"0ddd", x"0ddd", x"0ddd", x"0ddd", x"0ddd", x"0ddd", x"0ddd", x"0ddd", x"0ddd", x"0dde", x"0dde", x"0dde", x"0dde", x"0dde", x"0dde", x"0dde", x"0dde", x"0dde", x"0ddf", x"0ddf", x"0ddf", x"0ddf", x"0ddf", x"0ddf", x"0ddf", x"0ddf", x"0de0", x"0de0", x"0de0", x"0de0", x"0de0", x"0de0", x"0de0", x"0de0", x"0de0", x"0de1", x"0de1", x"0de1", x"0de1", x"0de1", x"0de1", x"0de1", x"0de1", x"0de1", x"0de2", x"0de2", x"0de2", x"0de2", x"0de2", x"0de2", x"0de2", x"0de2", x"0de2", x"0de3", x"0de3", x"0de3", x"0de3", x"0de3", x"0de3", x"0de3", x"0de3", x"0de4", x"0de4", x"0de4", x"0de4", x"0de4", x"0de4", x"0de4", x"0de4", x"0de4", x"0de5", x"0de5", x"0de5", x"0de5", x"0de5", x"0de5", x"0de5", x"0de5", x"0de5", x"0de6", x"0de6", x"0de6", x"0de6", x"0de6", x"0de6", x"0de6", x"0de6", x"0de6", x"0de7", x"0de7", x"0de7", x"0de7", x"0de7", x"0de7", x"0de7", x"0de7", x"0de8", x"0de8", x"0de8", x"0de8", x"0de8", x"0de8", x"0de8", x"0de8", x"0de8", x"0de9", x"0de9", x"0de9", x"0de9", x"0de9", x"0de9", x"0de9", x"0de9", x"0de9", x"0dea", x"0dea", x"0dea", x"0dea", x"0dea", x"0dea", x"0dea", x"0dea", x"0dea", x"0deb", x"0deb", x"0deb", x"0deb", x"0deb", x"0deb", x"0deb", x"0deb", x"0deb", x"0dec", x"0dec", x"0dec", x"0dec", x"0dec", x"0dec", x"0dec", x"0dec", x"0dec", x"0ded", x"0ded", x"0ded", x"0ded", x"0ded", x"0ded", x"0ded", x"0ded", x"0ded", x"0dee", x"0dee", x"0dee", x"0dee", x"0dee", x"0dee", x"0dee", x"0dee", x"0def", x"0def", x"0def", x"0def", x"0def", x"0def", x"0def", x"0def", x"0def", x"0df0", x"0df0", x"0df0", x"0df0", x"0df0", x"0df0", x"0df0", x"0df0", x"0df0", x"0df1", x"0df1", x"0df1", x"0df1", x"0df1", x"0df1", x"0df1", x"0df1", x"0df1", x"0df2", x"0df2", x"0df2", x"0df2", x"0df2", x"0df2", x"0df2", x"0df2", x"0df2", x"0df3", x"0df3", x"0df3", x"0df3", x"0df3", x"0df3", x"0df3", x"0df3", x"0df3", x"0df4", x"0df4", x"0df4", x"0df4", x"0df4", x"0df4", x"0df4", x"0df4", x"0df4", x"0df5", x"0df5", x"0df5", x"0df5", x"0df5", x"0df5", x"0df5", x"0df5", x"0df5", x"0df6", x"0df6", x"0df6", x"0df6", x"0df6", x"0df6", x"0df6", x"0df6", x"0df6", x"0df7", x"0df7", x"0df7", x"0df7", x"0df7", x"0df7", x"0df7", x"0df7", x"0df7", x"0df8", x"0df8", x"0df8", x"0df8", x"0df8", x"0df8", x"0df8", x"0df8", x"0df8", x"0df9", x"0df9", x"0df9", x"0df9", x"0df9", x"0df9", x"0df9", x"0df9", x"0df9", x"0dfa", x"0dfa", x"0dfa", x"0dfa", x"0dfa", x"0dfa", x"0dfa", x"0dfa", x"0dfa", x"0dfb", x"0dfb", x"0dfb", x"0dfb", x"0dfb", x"0dfb", x"0dfb", x"0dfb", x"0dfb", x"0dfc", x"0dfc", x"0dfc", x"0dfc", x"0dfc", x"0dfc", x"0dfc", x"0dfc", x"0dfc", x"0dfc", x"0dfd", x"0dfd", x"0dfd", x"0dfd", x"0dfd", x"0dfd", x"0dfd", x"0dfd", x"0dfd", x"0dfe", x"0dfe", x"0dfe", x"0dfe", x"0dfe", x"0dfe", x"0dfe", x"0dfe", x"0dfe", x"0dff", x"0dff", x"0dff", x"0dff", x"0dff", x"0dff", x"0dff", x"0dff", x"0dff", x"0e00", x"0e00", x"0e00", x"0e00", x"0e00", x"0e00", x"0e00", x"0e00", x"0e00", x"0e01", x"0e01", x"0e01", x"0e01", x"0e01", x"0e01", x"0e01", x"0e01", x"0e01", x"0e02", x"0e02", x"0e02", x"0e02", x"0e02", x"0e02", x"0e02", x"0e02", x"0e02", x"0e02", x"0e03", x"0e03", x"0e03", x"0e03", x"0e03", x"0e03", x"0e03", x"0e03", x"0e03", x"0e04", x"0e04", x"0e04", x"0e04", x"0e04", x"0e04", x"0e04", x"0e04", x"0e04", x"0e05", x"0e05", x"0e05", x"0e05", x"0e05", x"0e05", x"0e05", x"0e05", x"0e05", x"0e06", x"0e06", x"0e06", x"0e06", x"0e06", x"0e06", x"0e06", x"0e06", x"0e06", x"0e07", x"0e07", x"0e07", x"0e07", x"0e07", x"0e07", x"0e07", x"0e07", x"0e07", x"0e07", x"0e08", x"0e08", x"0e08", x"0e08", x"0e08", x"0e08", x"0e08", x"0e08", x"0e08", x"0e09", x"0e09", x"0e09", x"0e09", x"0e09", x"0e09", x"0e09", x"0e09", x"0e09", x"0e0a", x"0e0a", x"0e0a", x"0e0a", x"0e0a", x"0e0a", x"0e0a", x"0e0a", x"0e0a", x"0e0a", x"0e0b", x"0e0b", x"0e0b", x"0e0b", x"0e0b", x"0e0b", x"0e0b", x"0e0b", x"0e0b", x"0e0c", x"0e0c", x"0e0c", x"0e0c", x"0e0c", x"0e0c", x"0e0c", x"0e0c", x"0e0c", x"0e0d", x"0e0d", x"0e0d", x"0e0d", x"0e0d", x"0e0d", x"0e0d", x"0e0d", x"0e0d", x"0e0d", x"0e0e", x"0e0e", x"0e0e", x"0e0e", x"0e0e", x"0e0e", x"0e0e", x"0e0e", x"0e0e", x"0e0f", x"0e0f", x"0e0f", x"0e0f", x"0e0f", x"0e0f", x"0e0f", x"0e0f", x"0e0f", x"0e0f", x"0e10", x"0e10", x"0e10", x"0e10", x"0e10", x"0e10", x"0e10", x"0e10", x"0e10", x"0e11", x"0e11", x"0e11", x"0e11", x"0e11", x"0e11", x"0e11", x"0e11", x"0e11", x"0e12", x"0e12", x"0e12", x"0e12", x"0e12", x"0e12", x"0e12", x"0e12", x"0e12", x"0e12", x"0e13", x"0e13", x"0e13", x"0e13", x"0e13", x"0e13", x"0e13", x"0e13", x"0e13", x"0e14", x"0e14", x"0e14", x"0e14", x"0e14", x"0e14", x"0e14", x"0e14", x"0e14", x"0e14", x"0e15", x"0e15", x"0e15", x"0e15", x"0e15", x"0e15", x"0e15", x"0e15", x"0e15", x"0e16", x"0e16", x"0e16", x"0e16", x"0e16", x"0e16", x"0e16", x"0e16", x"0e16", x"0e16", x"0e17", x"0e17", x"0e17", x"0e17", x"0e17", x"0e17", x"0e17", x"0e17", x"0e17", x"0e18", x"0e18", x"0e18", x"0e18", x"0e18", x"0e18", x"0e18", x"0e18", x"0e18", x"0e18", x"0e19", x"0e19", x"0e19", x"0e19", x"0e19", x"0e19", x"0e19", x"0e19", x"0e19", x"0e1a", x"0e1a", x"0e1a", x"0e1a", x"0e1a", x"0e1a", x"0e1a", x"0e1a", x"0e1a", x"0e1a", x"0e1b", x"0e1b", x"0e1b", x"0e1b", x"0e1b", x"0e1b", x"0e1b", x"0e1b", x"0e1b", x"0e1b", x"0e1c", x"0e1c", x"0e1c", x"0e1c", x"0e1c", x"0e1c", x"0e1c", x"0e1c", x"0e1c", x"0e1d", x"0e1d", x"0e1d", x"0e1d", x"0e1d", x"0e1d", x"0e1d", x"0e1d", x"0e1d", x"0e1d", x"0e1e", x"0e1e", x"0e1e", x"0e1e", x"0e1e", x"0e1e", x"0e1e", x"0e1e", x"0e1e", x"0e1e", x"0e1f", x"0e1f", x"0e1f", x"0e1f", x"0e1f", x"0e1f", x"0e1f", x"0e1f", x"0e1f", x"0e20", x"0e20", x"0e20", x"0e20", x"0e20", x"0e20", x"0e20", x"0e20", x"0e20", x"0e20", x"0e21", x"0e21", x"0e21", x"0e21", x"0e21", x"0e21", x"0e21", x"0e21", x"0e21", x"0e21", x"0e22", x"0e22", x"0e22", x"0e22", x"0e22", x"0e22", x"0e22", x"0e22", x"0e22", x"0e23", x"0e23", x"0e23", x"0e23", x"0e23", x"0e23", x"0e23", x"0e23", x"0e23", x"0e23", x"0e24", x"0e24", x"0e24", x"0e24", x"0e24", x"0e24", x"0e24", x"0e24", x"0e24", x"0e24", x"0e25", x"0e25", x"0e25", x"0e25", x"0e25", x"0e25", x"0e25", x"0e25", x"0e25", x"0e25", x"0e26", x"0e26", x"0e26", x"0e26", x"0e26", x"0e26", x"0e26", x"0e26", x"0e26", x"0e27", x"0e27", x"0e27", x"0e27", x"0e27", x"0e27", x"0e27", x"0e27", x"0e27", x"0e27", x"0e28", x"0e28", x"0e28", x"0e28", x"0e28", x"0e28", x"0e28", x"0e28", x"0e28", x"0e28", x"0e29", x"0e29", x"0e29", x"0e29", x"0e29", x"0e29", x"0e29", x"0e29", x"0e29", x"0e29", x"0e2a", x"0e2a", x"0e2a", x"0e2a", x"0e2a", x"0e2a", x"0e2a", x"0e2a", x"0e2a", x"0e2a", x"0e2b", x"0e2b", x"0e2b", x"0e2b", x"0e2b", x"0e2b", x"0e2b", x"0e2b", x"0e2b", x"0e2b", x"0e2c", x"0e2c", x"0e2c", x"0e2c", x"0e2c", x"0e2c", x"0e2c", x"0e2c", x"0e2c", x"0e2c", x"0e2d", x"0e2d", x"0e2d", x"0e2d", x"0e2d", x"0e2d", x"0e2d", x"0e2d", x"0e2d", x"0e2d", x"0e2e", x"0e2e", x"0e2e", x"0e2e", x"0e2e", x"0e2e", x"0e2e", x"0e2e", x"0e2e", x"0e2e", x"0e2f", x"0e2f", x"0e2f", x"0e2f", x"0e2f", x"0e2f", x"0e2f", x"0e2f", x"0e2f", x"0e30", x"0e30", x"0e30", x"0e30", x"0e30", x"0e30", x"0e30", x"0e30", x"0e30", x"0e30", x"0e31", x"0e31", x"0e31", x"0e31", x"0e31", x"0e31", x"0e31", x"0e31", x"0e31", x"0e31", x"0e32", x"0e32", x"0e32", x"0e32", x"0e32", x"0e32", x"0e32", x"0e32", x"0e32", x"0e32", x"0e33", x"0e33", x"0e33", x"0e33", x"0e33", x"0e33", x"0e33", x"0e33", x"0e33", x"0e33", x"0e33", x"0e34", x"0e34", x"0e34", x"0e34", x"0e34", x"0e34", x"0e34", x"0e34", x"0e34", x"0e34", x"0e35", x"0e35", x"0e35", x"0e35", x"0e35", x"0e35", x"0e35", x"0e35", x"0e35", x"0e35", x"0e36", x"0e36", x"0e36", x"0e36", x"0e36", x"0e36", x"0e36", x"0e36", x"0e36", x"0e36", x"0e37", x"0e37", x"0e37", x"0e37", x"0e37", x"0e37", x"0e37", x"0e37", x"0e37", x"0e37", x"0e38", x"0e38", x"0e38", x"0e38", x"0e38", x"0e38", x"0e38", x"0e38", x"0e38", x"0e38", x"0e39", x"0e39", x"0e39", x"0e39", x"0e39", x"0e39", x"0e39", x"0e39", x"0e39", x"0e39", x"0e3a", x"0e3a", x"0e3a", x"0e3a", x"0e3a", x"0e3a", x"0e3a", x"0e3a", x"0e3a", x"0e3a", x"0e3b", x"0e3b", x"0e3b", x"0e3b", x"0e3b", x"0e3b", x"0e3b", x"0e3b", x"0e3b", x"0e3b", x"0e3b", x"0e3c", x"0e3c", x"0e3c", x"0e3c", x"0e3c", x"0e3c", x"0e3c", x"0e3c", x"0e3c", x"0e3c", x"0e3d", x"0e3d", x"0e3d", x"0e3d", x"0e3d", x"0e3d", x"0e3d", x"0e3d", x"0e3d", x"0e3d", x"0e3e", x"0e3e", x"0e3e", x"0e3e", x"0e3e", x"0e3e", x"0e3e", x"0e3e", x"0e3e", x"0e3e", x"0e3f", x"0e3f", x"0e3f", x"0e3f", x"0e3f", x"0e3f", x"0e3f", x"0e3f", x"0e3f", x"0e3f", x"0e3f", x"0e40", x"0e40", x"0e40", x"0e40", x"0e40", x"0e40", x"0e40", x"0e40", x"0e40", x"0e40", x"0e41", x"0e41", x"0e41", x"0e41", x"0e41", x"0e41", x"0e41", x"0e41", x"0e41", x"0e41", x"0e42", x"0e42", x"0e42", x"0e42", x"0e42", x"0e42", x"0e42", x"0e42", x"0e42", x"0e42", x"0e43", x"0e43", x"0e43", x"0e43", x"0e43", x"0e43", x"0e43", x"0e43", x"0e43", x"0e43", x"0e43", x"0e44", x"0e44", x"0e44", x"0e44", x"0e44", x"0e44", x"0e44", x"0e44", x"0e44", x"0e44", x"0e45", x"0e45", x"0e45", x"0e45", x"0e45", x"0e45", x"0e45", x"0e45", x"0e45", x"0e45", x"0e45", x"0e46", x"0e46", x"0e46", x"0e46", x"0e46", x"0e46", x"0e46", x"0e46", x"0e46", x"0e46", x"0e47", x"0e47", x"0e47", x"0e47", x"0e47", x"0e47", x"0e47", x"0e47", x"0e47", x"0e47", x"0e48", x"0e48", x"0e48", x"0e48", x"0e48", x"0e48", x"0e48", x"0e48", x"0e48", x"0e48", x"0e48", x"0e49", x"0e49", x"0e49", x"0e49", x"0e49", x"0e49", x"0e49", x"0e49", x"0e49", x"0e49", x"0e4a", x"0e4a", x"0e4a", x"0e4a", x"0e4a", x"0e4a", x"0e4a", x"0e4a", x"0e4a", x"0e4a", x"0e4a", x"0e4b", x"0e4b", x"0e4b", x"0e4b", x"0e4b", x"0e4b", x"0e4b", x"0e4b", x"0e4b", x"0e4b", x"0e4c", x"0e4c", x"0e4c", x"0e4c", x"0e4c", x"0e4c", x"0e4c", x"0e4c", x"0e4c", x"0e4c", x"0e4c", x"0e4d", x"0e4d", x"0e4d", x"0e4d", x"0e4d", x"0e4d", x"0e4d", x"0e4d", x"0e4d", x"0e4d", x"0e4d", x"0e4e", x"0e4e", x"0e4e", x"0e4e", x"0e4e", x"0e4e", x"0e4e", x"0e4e", x"0e4e", x"0e4e", x"0e4f", x"0e4f", x"0e4f", x"0e4f", x"0e4f", x"0e4f", x"0e4f", x"0e4f", x"0e4f", x"0e4f", x"0e4f", x"0e50", x"0e50", x"0e50", x"0e50", x"0e50", x"0e50", x"0e50", x"0e50", x"0e50", x"0e50", x"0e51", x"0e51", x"0e51", x"0e51", x"0e51", x"0e51", x"0e51", x"0e51", x"0e51", x"0e51", x"0e51", x"0e52", x"0e52", x"0e52", x"0e52", x"0e52", x"0e52", x"0e52", x"0e52", x"0e52", x"0e52", x"0e52", x"0e53", x"0e53", x"0e53", x"0e53", x"0e53", x"0e53", x"0e53", x"0e53", x"0e53", x"0e53", x"0e54", x"0e54", x"0e54", x"0e54", x"0e54", x"0e54", x"0e54", x"0e54", x"0e54", x"0e54", x"0e54", x"0e55", x"0e55", x"0e55", x"0e55", x"0e55", x"0e55", x"0e55", x"0e55", x"0e55", x"0e55", x"0e55", x"0e56", x"0e56", x"0e56", x"0e56", x"0e56", x"0e56", x"0e56", x"0e56", x"0e56", x"0e56", x"0e56", x"0e57", x"0e57", x"0e57", x"0e57", x"0e57", x"0e57", x"0e57", x"0e57", x"0e57", x"0e57", x"0e58", x"0e58", x"0e58", x"0e58", x"0e58", x"0e58", x"0e58", x"0e58", x"0e58", x"0e58", x"0e58", x"0e59", x"0e59", x"0e59", x"0e59", x"0e59", x"0e59", x"0e59", x"0e59", x"0e59", x"0e59", x"0e59", x"0e5a", x"0e5a", x"0e5a", x"0e5a", x"0e5a", x"0e5a", x"0e5a", x"0e5a", x"0e5a", x"0e5a", x"0e5a", x"0e5b", x"0e5b", x"0e5b", x"0e5b", x"0e5b", x"0e5b", x"0e5b", x"0e5b", x"0e5b", x"0e5b", x"0e5b", x"0e5c", x"0e5c", x"0e5c", x"0e5c", x"0e5c", x"0e5c", x"0e5c", x"0e5c", x"0e5c", x"0e5c", x"0e5c", x"0e5d", x"0e5d", x"0e5d", x"0e5d", x"0e5d", x"0e5d", x"0e5d", x"0e5d", x"0e5d", x"0e5d", x"0e5d", x"0e5e", x"0e5e", x"0e5e", x"0e5e", x"0e5e", x"0e5e", x"0e5e", x"0e5e", x"0e5e", x"0e5e", x"0e5e", x"0e5f", x"0e5f", x"0e5f", x"0e5f", x"0e5f", x"0e5f", x"0e5f", x"0e5f", x"0e5f", x"0e5f", x"0e5f", x"0e60", x"0e60", x"0e60", x"0e60", x"0e60", x"0e60", x"0e60", x"0e60", x"0e60", x"0e60", x"0e60", x"0e61", x"0e61", x"0e61", x"0e61", x"0e61", x"0e61", x"0e61", x"0e61", x"0e61", x"0e61", x"0e61", x"0e62", x"0e62", x"0e62", x"0e62", x"0e62", x"0e62", x"0e62", x"0e62", x"0e62", x"0e62", x"0e62", x"0e63", x"0e63", x"0e63", x"0e63", x"0e63", x"0e63", x"0e63", x"0e63", x"0e63", x"0e63", x"0e63", x"0e64", x"0e64", x"0e64", x"0e64", x"0e64", x"0e64", x"0e64", x"0e64", x"0e64", x"0e64", x"0e64", x"0e65", x"0e65", x"0e65", x"0e65", x"0e65", x"0e65", x"0e65", x"0e65", x"0e65", x"0e65", x"0e65", x"0e66", x"0e66", x"0e66", x"0e66", x"0e66", x"0e66", x"0e66", x"0e66", x"0e66", x"0e66", x"0e66", x"0e67", x"0e67", x"0e67", x"0e67", x"0e67", x"0e67", x"0e67", x"0e67", x"0e67", x"0e67", x"0e67", x"0e68", x"0e68", x"0e68", x"0e68", x"0e68", x"0e68", x"0e68", x"0e68", x"0e68", x"0e68", x"0e68", x"0e69", x"0e69", x"0e69", x"0e69", x"0e69", x"0e69", x"0e69", x"0e69", x"0e69", x"0e69", x"0e69", x"0e69", x"0e6a", x"0e6a", x"0e6a", x"0e6a", x"0e6a", x"0e6a", x"0e6a", x"0e6a", x"0e6a", x"0e6a", x"0e6a", x"0e6b", x"0e6b", x"0e6b", x"0e6b", x"0e6b", x"0e6b", x"0e6b", x"0e6b", x"0e6b", x"0e6b", x"0e6b", x"0e6c", x"0e6c", x"0e6c", x"0e6c", x"0e6c", x"0e6c", x"0e6c", x"0e6c", x"0e6c", x"0e6c", x"0e6c", x"0e6d", x"0e6d", x"0e6d", x"0e6d", x"0e6d", x"0e6d", x"0e6d", x"0e6d", x"0e6d", x"0e6d", x"0e6d", x"0e6d", x"0e6e", x"0e6e", x"0e6e", x"0e6e", x"0e6e", x"0e6e", x"0e6e", x"0e6e", x"0e6e", x"0e6e", x"0e6e", x"0e6f", x"0e6f", x"0e6f", x"0e6f", x"0e6f", x"0e6f", x"0e6f", x"0e6f", x"0e6f", x"0e6f", x"0e6f", x"0e70", x"0e70", x"0e70", x"0e70", x"0e70", x"0e70", x"0e70", x"0e70", x"0e70", x"0e70", x"0e70", x"0e70", x"0e71", x"0e71", x"0e71", x"0e71", x"0e71", x"0e71", x"0e71", x"0e71", x"0e71", x"0e71", x"0e71", x"0e72", x"0e72", x"0e72", x"0e72", x"0e72", x"0e72", x"0e72", x"0e72", x"0e72", x"0e72", x"0e72", x"0e72", x"0e73", x"0e73", x"0e73", x"0e73", x"0e73", x"0e73", x"0e73", x"0e73", x"0e73", x"0e73", x"0e73", x"0e74", x"0e74", x"0e74", x"0e74", x"0e74", x"0e74", x"0e74", x"0e74", x"0e74", x"0e74", x"0e74", x"0e74", x"0e75", x"0e75", x"0e75", x"0e75", x"0e75", x"0e75", x"0e75", x"0e75", x"0e75", x"0e75", x"0e75", x"0e76", x"0e76", x"0e76", x"0e76", x"0e76", x"0e76", x"0e76", x"0e76", x"0e76", x"0e76", x"0e76", x"0e76", x"0e77", x"0e77", x"0e77", x"0e77", x"0e77", x"0e77", x"0e77", x"0e77", x"0e77", x"0e77", x"0e77", x"0e78", x"0e78", x"0e78", x"0e78", x"0e78", x"0e78", x"0e78", x"0e78", x"0e78", x"0e78", x"0e78", x"0e78", x"0e79", x"0e79", x"0e79", x"0e79", x"0e79", x"0e79", x"0e79", x"0e79", x"0e79", x"0e79", x"0e79", x"0e7a", x"0e7a", x"0e7a", x"0e7a", x"0e7a", x"0e7a", x"0e7a", x"0e7a", x"0e7a", x"0e7a", x"0e7a", x"0e7a", x"0e7b", x"0e7b", x"0e7b", x"0e7b", x"0e7b", x"0e7b", x"0e7b", x"0e7b", x"0e7b", x"0e7b", x"0e7b", x"0e7b", x"0e7c", x"0e7c", x"0e7c", x"0e7c", x"0e7c", x"0e7c", x"0e7c", x"0e7c", x"0e7c", x"0e7c", x"0e7c", x"0e7d", x"0e7d", x"0e7d", x"0e7d", x"0e7d", x"0e7d", x"0e7d", x"0e7d", x"0e7d", x"0e7d", x"0e7d", x"0e7d", x"0e7e", x"0e7e", x"0e7e", x"0e7e", x"0e7e", x"0e7e", x"0e7e", x"0e7e", x"0e7e", x"0e7e", x"0e7e", x"0e7e", x"0e7f", x"0e7f", x"0e7f", x"0e7f", x"0e7f", x"0e7f", x"0e7f", x"0e7f", x"0e7f", x"0e7f", x"0e7f", x"0e7f", x"0e80", x"0e80", x"0e80", x"0e80", x"0e80", x"0e80", x"0e80", x"0e80", x"0e80", x"0e80", x"0e80", x"0e80", x"0e81", x"0e81", x"0e81", x"0e81", x"0e81", x"0e81", x"0e81", x"0e81", x"0e81", x"0e81", x"0e81", x"0e82", x"0e82", x"0e82", x"0e82", x"0e82", x"0e82", x"0e82", x"0e82", x"0e82", x"0e82", x"0e82", x"0e82", x"0e83", x"0e83", x"0e83", x"0e83", x"0e83", x"0e83", x"0e83", x"0e83", x"0e83", x"0e83", x"0e83", x"0e83", x"0e84", x"0e84", x"0e84", x"0e84", x"0e84", x"0e84", x"0e84", x"0e84", x"0e84", x"0e84", x"0e84", x"0e84", x"0e85", x"0e85", x"0e85", x"0e85", x"0e85", x"0e85", x"0e85", x"0e85", x"0e85", x"0e85", x"0e85", x"0e85", x"0e86", x"0e86", x"0e86", x"0e86", x"0e86", x"0e86", x"0e86", x"0e86", x"0e86", x"0e86", x"0e86", x"0e86", x"0e87", x"0e87", x"0e87", x"0e87", x"0e87", x"0e87", x"0e87", x"0e87", x"0e87", x"0e87", x"0e87", x"0e87", x"0e88", x"0e88", x"0e88", x"0e88", x"0e88", x"0e88", x"0e88", x"0e88", x"0e88", x"0e88", x"0e88", x"0e88", x"0e89", x"0e89", x"0e89", x"0e89", x"0e89", x"0e89", x"0e89", x"0e89", x"0e89", x"0e89", x"0e89", x"0e89", x"0e8a", x"0e8a", x"0e8a", x"0e8a", x"0e8a", x"0e8a", x"0e8a", x"0e8a", x"0e8a", x"0e8a", x"0e8a", x"0e8a", x"0e8b", x"0e8b", x"0e8b", x"0e8b", x"0e8b", x"0e8b", x"0e8b", x"0e8b", x"0e8b", x"0e8b", x"0e8b", x"0e8b", x"0e8c", x"0e8c", x"0e8c", x"0e8c", x"0e8c", x"0e8c", x"0e8c", x"0e8c", x"0e8c", x"0e8c", x"0e8c", x"0e8c", x"0e8d", x"0e8d", x"0e8d", x"0e8d", x"0e8d", x"0e8d", x"0e8d", x"0e8d", x"0e8d", x"0e8d", x"0e8d", x"0e8d", x"0e8d", x"0e8e", x"0e8e", x"0e8e", x"0e8e", x"0e8e", x"0e8e", x"0e8e", x"0e8e", x"0e8e", x"0e8e", x"0e8e", x"0e8e", x"0e8f", x"0e8f", x"0e8f", x"0e8f", x"0e8f", x"0e8f", x"0e8f", x"0e8f", x"0e8f", x"0e8f", x"0e8f", x"0e8f", x"0e90", x"0e90", x"0e90", x"0e90", x"0e90", x"0e90", x"0e90", x"0e90", x"0e90", x"0e90", x"0e90", x"0e90", x"0e91", x"0e91", x"0e91", x"0e91", x"0e91", x"0e91", x"0e91", x"0e91", x"0e91", x"0e91", x"0e91", x"0e91", x"0e91", x"0e92", x"0e92", x"0e92", x"0e92", x"0e92", x"0e92", x"0e92", x"0e92", x"0e92", x"0e92", x"0e92", x"0e92", x"0e93", x"0e93", x"0e93", x"0e93", x"0e93", x"0e93", x"0e93", x"0e93", x"0e93", x"0e93", x"0e93", x"0e93", x"0e94", x"0e94", x"0e94", x"0e94", x"0e94", x"0e94", x"0e94", x"0e94", x"0e94", x"0e94", x"0e94", x"0e94", x"0e94", x"0e95", x"0e95", x"0e95", x"0e95", x"0e95", x"0e95", x"0e95", x"0e95", x"0e95", x"0e95", x"0e95", x"0e95", x"0e96", x"0e96", x"0e96", x"0e96", x"0e96", x"0e96", x"0e96", x"0e96", x"0e96", x"0e96", x"0e96", x"0e96", x"0e96", x"0e97", x"0e97", x"0e97", x"0e97", x"0e97", x"0e97", x"0e97", x"0e97", x"0e97", x"0e97", x"0e97", x"0e97", x"0e98", x"0e98", x"0e98", x"0e98", x"0e98", x"0e98", x"0e98", x"0e98", x"0e98", x"0e98", x"0e98", x"0e98", x"0e98", x"0e99", x"0e99", x"0e99", x"0e99", x"0e99", x"0e99", x"0e99", x"0e99", x"0e99", x"0e99", x"0e99", x"0e99", x"0e9a", x"0e9a", x"0e9a", x"0e9a", x"0e9a", x"0e9a", x"0e9a", x"0e9a", x"0e9a", x"0e9a", x"0e9a", x"0e9a", x"0e9a", x"0e9b", x"0e9b", x"0e9b", x"0e9b", x"0e9b", x"0e9b", x"0e9b", x"0e9b", x"0e9b", x"0e9b", x"0e9b", x"0e9b", x"0e9c", x"0e9c", x"0e9c", x"0e9c", x"0e9c", x"0e9c", x"0e9c", x"0e9c", x"0e9c", x"0e9c", x"0e9c", x"0e9c", x"0e9c", x"0e9d", x"0e9d", x"0e9d", x"0e9d", x"0e9d", x"0e9d", x"0e9d", x"0e9d", x"0e9d", x"0e9d", x"0e9d", x"0e9d", x"0e9d", x"0e9e", x"0e9e", x"0e9e", x"0e9e", x"0e9e", x"0e9e", x"0e9e", x"0e9e", x"0e9e", x"0e9e", x"0e9e", x"0e9e", x"0e9f", x"0e9f", x"0e9f", x"0e9f", x"0e9f", x"0e9f", x"0e9f", x"0e9f", x"0e9f", x"0e9f", x"0e9f", x"0e9f", x"0e9f", x"0ea0", x"0ea0", x"0ea0", x"0ea0", x"0ea0", x"0ea0", x"0ea0", x"0ea0", x"0ea0", x"0ea0", x"0ea0", x"0ea0", x"0ea0", x"0ea1", x"0ea1", x"0ea1", x"0ea1", x"0ea1", x"0ea1", x"0ea1", x"0ea1", x"0ea1", x"0ea1", x"0ea1", x"0ea1", x"0ea1", x"0ea2", x"0ea2", x"0ea2", x"0ea2", x"0ea2", x"0ea2", x"0ea2", x"0ea2", x"0ea2", x"0ea2", x"0ea2", x"0ea2", x"0ea2", x"0ea3", x"0ea3", x"0ea3", x"0ea3", x"0ea3", x"0ea3", x"0ea3", x"0ea3", x"0ea3", x"0ea3", x"0ea3", x"0ea3", x"0ea3", x"0ea4", x"0ea4", x"0ea4", x"0ea4", x"0ea4", x"0ea4", x"0ea4", x"0ea4", x"0ea4", x"0ea4", x"0ea4", x"0ea4", x"0ea5", x"0ea5", x"0ea5", x"0ea5", x"0ea5", x"0ea5", x"0ea5", x"0ea5", x"0ea5", x"0ea5", x"0ea5", x"0ea5", x"0ea5", x"0ea6", x"0ea6", x"0ea6", x"0ea6", x"0ea6", x"0ea6", x"0ea6", x"0ea6", x"0ea6", x"0ea6", x"0ea6", x"0ea6", x"0ea6", x"0ea7", x"0ea7", x"0ea7", x"0ea7", x"0ea7", x"0ea7", x"0ea7", x"0ea7", x"0ea7", x"0ea7", x"0ea7", x"0ea7", x"0ea7", x"0ea8", x"0ea8", x"0ea8", x"0ea8", x"0ea8", x"0ea8", x"0ea8", x"0ea8", x"0ea8", x"0ea8", x"0ea8", x"0ea8", x"0ea8", x"0ea9", x"0ea9", x"0ea9", x"0ea9", x"0ea9", x"0ea9", x"0ea9", x"0ea9", x"0ea9", x"0ea9", x"0ea9", x"0ea9", x"0ea9", x"0ea9", x"0eaa", x"0eaa", x"0eaa", x"0eaa", x"0eaa", x"0eaa", x"0eaa", x"0eaa", x"0eaa", x"0eaa", x"0eaa", x"0eaa", x"0eaa", x"0eab", x"0eab", x"0eab", x"0eab", x"0eab", x"0eab", x"0eab", x"0eab", x"0eab", x"0eab", x"0eab", x"0eab", x"0eab", x"0eac", x"0eac", x"0eac", x"0eac", x"0eac", x"0eac", x"0eac", x"0eac", x"0eac", x"0eac", x"0eac", x"0eac", x"0eac", x"0ead", x"0ead", x"0ead", x"0ead", x"0ead", x"0ead", x"0ead", x"0ead", x"0ead", x"0ead", x"0ead", x"0ead", x"0ead", x"0eae", x"0eae", x"0eae", x"0eae", x"0eae", x"0eae", x"0eae", x"0eae", x"0eae", x"0eae", x"0eae", x"0eae", x"0eae", x"0eae", x"0eaf", x"0eaf", x"0eaf", x"0eaf", x"0eaf", x"0eaf", x"0eaf", x"0eaf", x"0eaf", x"0eaf", x"0eaf", x"0eaf", x"0eaf", x"0eb0", x"0eb0", x"0eb0", x"0eb0", x"0eb0", x"0eb0", x"0eb0", x"0eb0", x"0eb0", x"0eb0", x"0eb0", x"0eb0", x"0eb0", x"0eb1", x"0eb1", x"0eb1", x"0eb1", x"0eb1", x"0eb1", x"0eb1", x"0eb1", x"0eb1", x"0eb1", x"0eb1", x"0eb1", x"0eb1", x"0eb1", x"0eb2", x"0eb2", x"0eb2", x"0eb2", x"0eb2", x"0eb2", x"0eb2", x"0eb2", x"0eb2", x"0eb2", x"0eb2", x"0eb2", x"0eb2", x"0eb3", x"0eb3", x"0eb3", x"0eb3", x"0eb3", x"0eb3", x"0eb3", x"0eb3", x"0eb3", x"0eb3", x"0eb3", x"0eb3", x"0eb3", x"0eb4", x"0eb4", x"0eb4", x"0eb4", x"0eb4", x"0eb4", x"0eb4", x"0eb4", x"0eb4", x"0eb4", x"0eb4", x"0eb4", x"0eb4", x"0eb4", x"0eb5", x"0eb5", x"0eb5", x"0eb5", x"0eb5", x"0eb5", x"0eb5", x"0eb5", x"0eb5", x"0eb5", x"0eb5", x"0eb5", x"0eb5", x"0eb6", x"0eb6", x"0eb6", x"0eb6", x"0eb6", x"0eb6", x"0eb6", x"0eb6", x"0eb6", x"0eb6", x"0eb6", x"0eb6", x"0eb6", x"0eb6", x"0eb7", x"0eb7", x"0eb7", x"0eb7", x"0eb7", x"0eb7", x"0eb7", x"0eb7", x"0eb7", x"0eb7", x"0eb7", x"0eb7", x"0eb7", x"0eb7", x"0eb8", x"0eb8", x"0eb8", x"0eb8", x"0eb8", x"0eb8", x"0eb8", x"0eb8", x"0eb8", x"0eb8", x"0eb8", x"0eb8", x"0eb8", x"0eb9", x"0eb9", x"0eb9", x"0eb9", x"0eb9", x"0eb9", x"0eb9", x"0eb9", x"0eb9", x"0eb9", x"0eb9", x"0eb9", x"0eb9", x"0eb9", x"0eba", x"0eba", x"0eba", x"0eba", x"0eba", x"0eba", x"0eba", x"0eba", x"0eba", x"0eba", x"0eba", x"0eba", x"0eba", x"0eba", x"0ebb", x"0ebb", x"0ebb", x"0ebb", x"0ebb", x"0ebb", x"0ebb", x"0ebb", x"0ebb", x"0ebb", x"0ebb", x"0ebb", x"0ebb", x"0ebc", x"0ebc", x"0ebc", x"0ebc", x"0ebc", x"0ebc", x"0ebc", x"0ebc", x"0ebc", x"0ebc", x"0ebc", x"0ebc", x"0ebc", x"0ebc", x"0ebd", x"0ebd", x"0ebd", x"0ebd", x"0ebd", x"0ebd", x"0ebd", x"0ebd", x"0ebd", x"0ebd", x"0ebd", x"0ebd", x"0ebd", x"0ebd", x"0ebe", x"0ebe", x"0ebe", x"0ebe", x"0ebe", x"0ebe", x"0ebe", x"0ebe", x"0ebe", x"0ebe", x"0ebe", x"0ebe", x"0ebe", x"0ebe", x"0ebf", x"0ebf", x"0ebf", x"0ebf", x"0ebf", x"0ebf", x"0ebf", x"0ebf", x"0ebf", x"0ebf", x"0ebf", x"0ebf", x"0ebf", x"0ebf", x"0ec0", x"0ec0", x"0ec0", x"0ec0", x"0ec0", x"0ec0", x"0ec0", x"0ec0", x"0ec0", x"0ec0", x"0ec0", x"0ec0", x"0ec0", x"0ec0", x"0ec1", x"0ec1", x"0ec1", x"0ec1", x"0ec1", x"0ec1", x"0ec1", x"0ec1", x"0ec1", x"0ec1", x"0ec1", x"0ec1", x"0ec1", x"0ec1", x"0ec2", x"0ec2", x"0ec2", x"0ec2", x"0ec2", x"0ec2", x"0ec2", x"0ec2", x"0ec2", x"0ec2", x"0ec2", x"0ec2", x"0ec2", x"0ec2", x"0ec3", x"0ec3", x"0ec3", x"0ec3", x"0ec3", x"0ec3", x"0ec3", x"0ec3", x"0ec3", x"0ec3", x"0ec3", x"0ec3", x"0ec3", x"0ec3", x"0ec4", x"0ec4", x"0ec4", x"0ec4", x"0ec4", x"0ec4", x"0ec4", x"0ec4", x"0ec4", x"0ec4", x"0ec4", x"0ec4", x"0ec4", x"0ec4", x"0ec5", x"0ec5", x"0ec5", x"0ec5", x"0ec5", x"0ec5", x"0ec5", x"0ec5", x"0ec5", x"0ec5", x"0ec5", x"0ec5", x"0ec5", x"0ec5", x"0ec6", x"0ec6", x"0ec6", x"0ec6", x"0ec6", x"0ec6", x"0ec6", x"0ec6", x"0ec6", x"0ec6", x"0ec6", x"0ec6", x"0ec6", x"0ec6", x"0ec7", x"0ec7", x"0ec7", x"0ec7", x"0ec7", x"0ec7", x"0ec7", x"0ec7", x"0ec7", x"0ec7", x"0ec7", x"0ec7", x"0ec7", x"0ec7", x"0ec8", x"0ec8", x"0ec8", x"0ec8", x"0ec8", x"0ec8", x"0ec8", x"0ec8", x"0ec8", x"0ec8", x"0ec8", x"0ec8", x"0ec8", x"0ec8", x"0ec8", x"0ec9", x"0ec9", x"0ec9", x"0ec9", x"0ec9", x"0ec9", x"0ec9", x"0ec9", x"0ec9", x"0ec9", x"0ec9", x"0ec9", x"0ec9", x"0ec9", x"0eca", x"0eca", x"0eca", x"0eca", x"0eca", x"0eca", x"0eca", x"0eca", x"0eca", x"0eca", x"0eca", x"0eca", x"0eca", x"0eca", x"0ecb", x"0ecb", x"0ecb", x"0ecb", x"0ecb", x"0ecb", x"0ecb", x"0ecb", x"0ecb", x"0ecb", x"0ecb", x"0ecb", x"0ecb", x"0ecb", x"0ecb", x"0ecc", x"0ecc", x"0ecc", x"0ecc", x"0ecc", x"0ecc", x"0ecc", x"0ecc", x"0ecc", x"0ecc", x"0ecc", x"0ecc", x"0ecc", x"0ecc", x"0ecd", x"0ecd", x"0ecd", x"0ecd", x"0ecd", x"0ecd", x"0ecd", x"0ecd", x"0ecd", x"0ecd", x"0ecd", x"0ecd", x"0ecd", x"0ecd", x"0ecd", x"0ece", x"0ece", x"0ece", x"0ece", x"0ece", x"0ece", x"0ece", x"0ece", x"0ece", x"0ece", x"0ece", x"0ece", x"0ece", x"0ece", x"0ecf", x"0ecf", x"0ecf", x"0ecf", x"0ecf", x"0ecf", x"0ecf", x"0ecf", x"0ecf", x"0ecf", x"0ecf", x"0ecf", x"0ecf", x"0ecf", x"0ecf", x"0ed0", x"0ed0", x"0ed0", x"0ed0", x"0ed0", x"0ed0", x"0ed0", x"0ed0", x"0ed0", x"0ed0", x"0ed0", x"0ed0", x"0ed0", x"0ed0", x"0ed1", x"0ed1", x"0ed1", x"0ed1", x"0ed1", x"0ed1", x"0ed1", x"0ed1", x"0ed1", x"0ed1", x"0ed1", x"0ed1", x"0ed1", x"0ed1", x"0ed1", x"0ed2", x"0ed2", x"0ed2", x"0ed2", x"0ed2", x"0ed2", x"0ed2", x"0ed2", x"0ed2", x"0ed2", x"0ed2", x"0ed2", x"0ed2", x"0ed2", x"0ed2", x"0ed3", x"0ed3", x"0ed3", x"0ed3", x"0ed3", x"0ed3", x"0ed3", x"0ed3", x"0ed3", x"0ed3", x"0ed3", x"0ed3", x"0ed3", x"0ed3", x"0ed4", x"0ed4", x"0ed4", x"0ed4", x"0ed4", x"0ed4", x"0ed4", x"0ed4", x"0ed4", x"0ed4", x"0ed4", x"0ed4", x"0ed4", x"0ed4", x"0ed4", x"0ed5", x"0ed5", x"0ed5", x"0ed5", x"0ed5", x"0ed5", x"0ed5", x"0ed5", x"0ed5", x"0ed5", x"0ed5", x"0ed5", x"0ed5", x"0ed5", x"0ed5", x"0ed6", x"0ed6", x"0ed6", x"0ed6", x"0ed6", x"0ed6", x"0ed6", x"0ed6", x"0ed6", x"0ed6", x"0ed6", x"0ed6", x"0ed6", x"0ed6", x"0ed6", x"0ed7", x"0ed7", x"0ed7", x"0ed7", x"0ed7", x"0ed7", x"0ed7", x"0ed7", x"0ed7", x"0ed7", x"0ed7", x"0ed7", x"0ed7", x"0ed7", x"0ed7", x"0ed8", x"0ed8", x"0ed8", x"0ed8", x"0ed8", x"0ed8", x"0ed8", x"0ed8", x"0ed8", x"0ed8", x"0ed8", x"0ed8", x"0ed8", x"0ed8", x"0ed8", x"0ed9", x"0ed9", x"0ed9", x"0ed9", x"0ed9", x"0ed9", x"0ed9", x"0ed9", x"0ed9", x"0ed9", x"0ed9", x"0ed9", x"0ed9", x"0ed9", x"0ed9", x"0eda", x"0eda", x"0eda", x"0eda", x"0eda", x"0eda", x"0eda", x"0eda", x"0eda", x"0eda", x"0eda", x"0eda", x"0eda", x"0eda", x"0eda", x"0edb", x"0edb", x"0edb", x"0edb", x"0edb", x"0edb", x"0edb", x"0edb", x"0edb", x"0edb", x"0edb", x"0edb", x"0edb", x"0edb", x"0edb", x"0edc", x"0edc", x"0edc", x"0edc", x"0edc", x"0edc", x"0edc", x"0edc", x"0edc", x"0edc", x"0edc", x"0edc", x"0edc", x"0edc", x"0edc", x"0edd", x"0edd", x"0edd", x"0edd", x"0edd", x"0edd", x"0edd", x"0edd", x"0edd", x"0edd", x"0edd", x"0edd", x"0edd", x"0edd", x"0edd", x"0edd", x"0ede", x"0ede", x"0ede", x"0ede", x"0ede", x"0ede", x"0ede", x"0ede", x"0ede", x"0ede", x"0ede", x"0ede", x"0ede", x"0ede", x"0ede", x"0edf", x"0edf", x"0edf", x"0edf", x"0edf", x"0edf", x"0edf", x"0edf", x"0edf", x"0edf", x"0edf", x"0edf", x"0edf", x"0edf", x"0edf", x"0ee0", x"0ee0", x"0ee0", x"0ee0", x"0ee0", x"0ee0", x"0ee0", x"0ee0", x"0ee0", x"0ee0", x"0ee0", x"0ee0", x"0ee0", x"0ee0", x"0ee0", x"0ee0", x"0ee1", x"0ee1", x"0ee1", x"0ee1", x"0ee1", x"0ee1", x"0ee1", x"0ee1", x"0ee1", x"0ee1", x"0ee1", x"0ee1", x"0ee1", x"0ee1", x"0ee1", x"0ee2", x"0ee2", x"0ee2", x"0ee2", x"0ee2", x"0ee2", x"0ee2", x"0ee2", x"0ee2", x"0ee2", x"0ee2", x"0ee2", x"0ee2", x"0ee2", x"0ee2", x"0ee3", x"0ee3", x"0ee3", x"0ee3", x"0ee3", x"0ee3", x"0ee3", x"0ee3", x"0ee3", x"0ee3", x"0ee3", x"0ee3", x"0ee3", x"0ee3", x"0ee3", x"0ee3", x"0ee4", x"0ee4", x"0ee4", x"0ee4", x"0ee4", x"0ee4", x"0ee4", x"0ee4", x"0ee4", x"0ee4", x"0ee4", x"0ee4", x"0ee4", x"0ee4", x"0ee4", x"0ee4", x"0ee5", x"0ee5", x"0ee5", x"0ee5", x"0ee5", x"0ee5", x"0ee5", x"0ee5", x"0ee5", x"0ee5", x"0ee5", x"0ee5", x"0ee5", x"0ee5", x"0ee5", x"0ee6", x"0ee6", x"0ee6", x"0ee6", x"0ee6", x"0ee6", x"0ee6", x"0ee6", x"0ee6", x"0ee6", x"0ee6", x"0ee6", x"0ee6", x"0ee6", x"0ee6", x"0ee6", x"0ee7", x"0ee7", x"0ee7", x"0ee7", x"0ee7", x"0ee7", x"0ee7", x"0ee7", x"0ee7", x"0ee7", x"0ee7", x"0ee7", x"0ee7", x"0ee7", x"0ee7", x"0ee7", x"0ee8", x"0ee8", x"0ee8", x"0ee8", x"0ee8", x"0ee8", x"0ee8", x"0ee8", x"0ee8", x"0ee8", x"0ee8", x"0ee8", x"0ee8", x"0ee8", x"0ee8", x"0ee9", x"0ee9", x"0ee9", x"0ee9", x"0ee9", x"0ee9", x"0ee9", x"0ee9", x"0ee9", x"0ee9", x"0ee9", x"0ee9", x"0ee9", x"0ee9", x"0ee9", x"0ee9", x"0eea", x"0eea", x"0eea", x"0eea", x"0eea", x"0eea", x"0eea", x"0eea", x"0eea", x"0eea", x"0eea", x"0eea", x"0eea", x"0eea", x"0eea", x"0eea", x"0eeb", x"0eeb", x"0eeb", x"0eeb", x"0eeb", x"0eeb", x"0eeb", x"0eeb", x"0eeb", x"0eeb", x"0eeb", x"0eeb", x"0eeb", x"0eeb", x"0eeb", x"0eeb", x"0eec", x"0eec", x"0eec", x"0eec", x"0eec", x"0eec", x"0eec", x"0eec", x"0eec", x"0eec", x"0eec", x"0eec", x"0eec", x"0eec", x"0eec", x"0eec", x"0eed", x"0eed", x"0eed", x"0eed", x"0eed", x"0eed", x"0eed", x"0eed", x"0eed", x"0eed", x"0eed", x"0eed", x"0eed", x"0eed", x"0eed", x"0eed", x"0eee", x"0eee", x"0eee", x"0eee", x"0eee", x"0eee", x"0eee", x"0eee", x"0eee", x"0eee", x"0eee", x"0eee", x"0eee", x"0eee", x"0eee", x"0eee", x"0eef", x"0eef", x"0eef", x"0eef", x"0eef", x"0eef", x"0eef", x"0eef", x"0eef", x"0eef", x"0eef", x"0eef", x"0eef", x"0eef", x"0eef", x"0eef", x"0ef0", x"0ef0", x"0ef0", x"0ef0", x"0ef0", x"0ef0", x"0ef0", x"0ef0", x"0ef0", x"0ef0", x"0ef0", x"0ef0", x"0ef0", x"0ef0", x"0ef0", x"0ef0", x"0ef0", x"0ef1", x"0ef1", x"0ef1", x"0ef1", x"0ef1", x"0ef1", x"0ef1", x"0ef1", x"0ef1", x"0ef1", x"0ef1", x"0ef1", x"0ef1", x"0ef1", x"0ef1", x"0ef1", x"0ef2", x"0ef2", x"0ef2", x"0ef2", x"0ef2", x"0ef2", x"0ef2", x"0ef2", x"0ef2", x"0ef2", x"0ef2", x"0ef2", x"0ef2", x"0ef2", x"0ef2", x"0ef2", x"0ef3", x"0ef3", x"0ef3", x"0ef3", x"0ef3", x"0ef3", x"0ef3", x"0ef3", x"0ef3", x"0ef3", x"0ef3", x"0ef3", x"0ef3", x"0ef3", x"0ef3", x"0ef3", x"0ef3", x"0ef4", x"0ef4", x"0ef4", x"0ef4", x"0ef4", x"0ef4", x"0ef4", x"0ef4", x"0ef4", x"0ef4", x"0ef4", x"0ef4", x"0ef4", x"0ef4", x"0ef4", x"0ef4", x"0ef5", x"0ef5", x"0ef5", x"0ef5", x"0ef5", x"0ef5", x"0ef5", x"0ef5", x"0ef5", x"0ef5", x"0ef5", x"0ef5", x"0ef5", x"0ef5", x"0ef5", x"0ef5", x"0ef6", x"0ef6", x"0ef6", x"0ef6", x"0ef6", x"0ef6", x"0ef6", x"0ef6", x"0ef6", x"0ef6", x"0ef6", x"0ef6", x"0ef6", x"0ef6", x"0ef6", x"0ef6", x"0ef6", x"0ef7", x"0ef7", x"0ef7", x"0ef7", x"0ef7", x"0ef7", x"0ef7", x"0ef7", x"0ef7", x"0ef7", x"0ef7", x"0ef7", x"0ef7", x"0ef7", x"0ef7", x"0ef7", x"0ef7", x"0ef8", x"0ef8", x"0ef8", x"0ef8", x"0ef8", x"0ef8", x"0ef8", x"0ef8", x"0ef8", x"0ef8", x"0ef8", x"0ef8", x"0ef8", x"0ef8", x"0ef8", x"0ef8", x"0ef9", x"0ef9", x"0ef9", x"0ef9", x"0ef9", x"0ef9", x"0ef9", x"0ef9", x"0ef9", x"0ef9", x"0ef9", x"0ef9", x"0ef9", x"0ef9", x"0ef9", x"0ef9", x"0ef9", x"0efa", x"0efa", x"0efa", x"0efa", x"0efa", x"0efa", x"0efa", x"0efa", x"0efa", x"0efa", x"0efa", x"0efa", x"0efa", x"0efa", x"0efa", x"0efa", x"0efa", x"0efb", x"0efb", x"0efb", x"0efb", x"0efb", x"0efb", x"0efb", x"0efb", x"0efb", x"0efb", x"0efb", x"0efb", x"0efb", x"0efb", x"0efb", x"0efb", x"0efb", x"0efc", x"0efc", x"0efc", x"0efc", x"0efc", x"0efc", x"0efc", x"0efc", x"0efc", x"0efc", x"0efc", x"0efc", x"0efc", x"0efc", x"0efc", x"0efc", x"0efc", x"0efd", x"0efd", x"0efd", x"0efd", x"0efd", x"0efd", x"0efd", x"0efd", x"0efd", x"0efd", x"0efd", x"0efd", x"0efd", x"0efd", x"0efd", x"0efd", x"0efd", x"0efe", x"0efe", x"0efe", x"0efe", x"0efe", x"0efe", x"0efe", x"0efe", x"0efe", x"0efe", x"0efe", x"0efe", x"0efe", x"0efe", x"0efe", x"0efe", x"0efe", x"0eff", x"0eff", x"0eff", x"0eff", x"0eff", x"0eff", x"0eff", x"0eff", x"0eff", x"0eff", x"0eff", x"0eff", x"0eff", x"0eff", x"0eff", x"0eff", x"0eff", x"0f00", x"0f00", x"0f00", x"0f00", x"0f00", x"0f00", x"0f00", x"0f00", x"0f00", x"0f00", x"0f00", x"0f00", x"0f00", x"0f00", x"0f00", x"0f00", x"0f00", x"0f01", x"0f01", x"0f01", x"0f01", x"0f01", x"0f01", x"0f01", x"0f01", x"0f01", x"0f01", x"0f01", x"0f01", x"0f01", x"0f01", x"0f01", x"0f01", x"0f01", x"0f02", x"0f02", x"0f02", x"0f02", x"0f02", x"0f02", x"0f02", x"0f02", x"0f02", x"0f02", x"0f02", x"0f02", x"0f02", x"0f02", x"0f02", x"0f02", x"0f02", x"0f03", x"0f03", x"0f03", x"0f03", x"0f03", x"0f03", x"0f03", x"0f03", x"0f03", x"0f03", x"0f03", x"0f03", x"0f03", x"0f03", x"0f03", x"0f03", x"0f03", x"0f03", x"0f04", x"0f04", x"0f04", x"0f04", x"0f04", x"0f04", x"0f04", x"0f04", x"0f04", x"0f04", x"0f04", x"0f04", x"0f04", x"0f04", x"0f04", x"0f04", x"0f04", x"0f05", x"0f05", x"0f05", x"0f05", x"0f05", x"0f05", x"0f05", x"0f05", x"0f05", x"0f05", x"0f05", x"0f05", x"0f05", x"0f05", x"0f05", x"0f05", x"0f05", x"0f05", x"0f06", x"0f06", x"0f06", x"0f06", x"0f06", x"0f06", x"0f06", x"0f06", x"0f06", x"0f06", x"0f06", x"0f06", x"0f06", x"0f06", x"0f06", x"0f06", x"0f06", x"0f07", x"0f07", x"0f07", x"0f07", x"0f07", x"0f07", x"0f07", x"0f07", x"0f07", x"0f07", x"0f07", x"0f07", x"0f07", x"0f07", x"0f07", x"0f07", x"0f07", x"0f07", x"0f08", x"0f08", x"0f08", x"0f08", x"0f08", x"0f08", x"0f08", x"0f08", x"0f08", x"0f08", x"0f08", x"0f08", x"0f08", x"0f08", x"0f08", x"0f08", x"0f08", x"0f09", x"0f09", x"0f09", x"0f09", x"0f09", x"0f09", x"0f09", x"0f09", x"0f09", x"0f09", x"0f09", x"0f09", x"0f09", x"0f09", x"0f09", x"0f09", x"0f09", x"0f09", x"0f0a", x"0f0a", x"0f0a", x"0f0a", x"0f0a", x"0f0a", x"0f0a", x"0f0a", x"0f0a", x"0f0a", x"0f0a", x"0f0a", x"0f0a", x"0f0a", x"0f0a", x"0f0a", x"0f0a", x"0f0a", x"0f0b", x"0f0b", x"0f0b", x"0f0b", x"0f0b", x"0f0b", x"0f0b", x"0f0b", x"0f0b", x"0f0b", x"0f0b", x"0f0b", x"0f0b", x"0f0b", x"0f0b", x"0f0b", x"0f0b", x"0f0b", x"0f0c", x"0f0c", x"0f0c", x"0f0c", x"0f0c", x"0f0c", x"0f0c", x"0f0c", x"0f0c", x"0f0c", x"0f0c", x"0f0c", x"0f0c", x"0f0c", x"0f0c", x"0f0c", x"0f0c", x"0f0c", x"0f0d", x"0f0d", x"0f0d", x"0f0d", x"0f0d", x"0f0d", x"0f0d", x"0f0d", x"0f0d", x"0f0d", x"0f0d", x"0f0d", x"0f0d", x"0f0d", x"0f0d", x"0f0d", x"0f0d", x"0f0d", x"0f0e", x"0f0e", x"0f0e", x"0f0e", x"0f0e", x"0f0e", x"0f0e", x"0f0e", x"0f0e", x"0f0e", x"0f0e", x"0f0e", x"0f0e", x"0f0e", x"0f0e", x"0f0e", x"0f0e", x"0f0e", x"0f0f", x"0f0f", x"0f0f", x"0f0f", x"0f0f", x"0f0f", x"0f0f", x"0f0f", x"0f0f", x"0f0f", x"0f0f", x"0f0f", x"0f0f", x"0f0f", x"0f0f", x"0f0f", x"0f0f", x"0f0f", x"0f10", x"0f10", x"0f10", x"0f10", x"0f10", x"0f10", x"0f10", x"0f10", x"0f10", x"0f10", x"0f10", x"0f10", x"0f10", x"0f10", x"0f10", x"0f10", x"0f10", x"0f10", x"0f11", x"0f11", x"0f11", x"0f11", x"0f11", x"0f11", x"0f11", x"0f11", x"0f11", x"0f11", x"0f11", x"0f11", x"0f11", x"0f11", x"0f11", x"0f11", x"0f11", x"0f11", x"0f11", x"0f12", x"0f12", x"0f12", x"0f12", x"0f12", x"0f12", x"0f12", x"0f12", x"0f12", x"0f12", x"0f12", x"0f12", x"0f12", x"0f12", x"0f12", x"0f12", x"0f12", x"0f12", x"0f13", x"0f13", x"0f13", x"0f13", x"0f13", x"0f13", x"0f13", x"0f13", x"0f13", x"0f13", x"0f13", x"0f13", x"0f13", x"0f13", x"0f13", x"0f13", x"0f13", x"0f13", x"0f13", x"0f14", x"0f14", x"0f14", x"0f14", x"0f14", x"0f14", x"0f14", x"0f14", x"0f14", x"0f14", x"0f14", x"0f14", x"0f14", x"0f14", x"0f14", x"0f14", x"0f14", x"0f14", x"0f15", x"0f15", x"0f15", x"0f15", x"0f15", x"0f15", x"0f15", x"0f15", x"0f15", x"0f15", x"0f15", x"0f15", x"0f15", x"0f15", x"0f15", x"0f15", x"0f15", x"0f15", x"0f15", x"0f16", x"0f16", x"0f16", x"0f16", x"0f16", x"0f16", x"0f16", x"0f16", x"0f16", x"0f16", x"0f16", x"0f16", x"0f16", x"0f16", x"0f16", x"0f16", x"0f16", x"0f16", x"0f17", x"0f17", x"0f17", x"0f17", x"0f17", x"0f17", x"0f17", x"0f17", x"0f17", x"0f17", x"0f17", x"0f17", x"0f17", x"0f17", x"0f17", x"0f17", x"0f17", x"0f17", x"0f17", x"0f18", x"0f18", x"0f18", x"0f18", x"0f18", x"0f18", x"0f18", x"0f18", x"0f18", x"0f18", x"0f18", x"0f18", x"0f18", x"0f18", x"0f18", x"0f18", x"0f18", x"0f18", x"0f18", x"0f19", x"0f19", x"0f19", x"0f19", x"0f19", x"0f19", x"0f19", x"0f19", x"0f19", x"0f19", x"0f19", x"0f19", x"0f19", x"0f19", x"0f19", x"0f19", x"0f19", x"0f19", x"0f19", x"0f1a", x"0f1a", x"0f1a", x"0f1a", x"0f1a", x"0f1a", x"0f1a", x"0f1a", x"0f1a", x"0f1a", x"0f1a", x"0f1a", x"0f1a", x"0f1a", x"0f1a", x"0f1a", x"0f1a", x"0f1a", x"0f1a", x"0f1b", x"0f1b", x"0f1b", x"0f1b", x"0f1b", x"0f1b", x"0f1b", x"0f1b", x"0f1b", x"0f1b", x"0f1b", x"0f1b", x"0f1b", x"0f1b", x"0f1b", x"0f1b", x"0f1b", x"0f1b", x"0f1b", x"0f1c", x"0f1c", x"0f1c", x"0f1c", x"0f1c", x"0f1c", x"0f1c", x"0f1c", x"0f1c", x"0f1c", x"0f1c", x"0f1c", x"0f1c", x"0f1c", x"0f1c", x"0f1c", x"0f1c", x"0f1c", x"0f1c", x"0f1d", x"0f1d", x"0f1d", x"0f1d", x"0f1d", x"0f1d", x"0f1d", x"0f1d", x"0f1d", x"0f1d", x"0f1d", x"0f1d", x"0f1d", x"0f1d", x"0f1d", x"0f1d", x"0f1d", x"0f1d", x"0f1d", x"0f1e", x"0f1e", x"0f1e", x"0f1e", x"0f1e", x"0f1e", x"0f1e", x"0f1e", x"0f1e", x"0f1e", x"0f1e", x"0f1e", x"0f1e", x"0f1e", x"0f1e", x"0f1e", x"0f1e", x"0f1e", x"0f1e", x"0f1e", x"0f1f", x"0f1f", x"0f1f", x"0f1f", x"0f1f", x"0f1f", x"0f1f", x"0f1f", x"0f1f", x"0f1f", x"0f1f", x"0f1f", x"0f1f", x"0f1f", x"0f1f", x"0f1f", x"0f1f", x"0f1f", x"0f1f", x"0f20", x"0f20", x"0f20", x"0f20", x"0f20", x"0f20", x"0f20", x"0f20", x"0f20", x"0f20", x"0f20", x"0f20", x"0f20", x"0f20", x"0f20", x"0f20", x"0f20", x"0f20", x"0f20", x"0f21", x"0f21", x"0f21", x"0f21", x"0f21", x"0f21", x"0f21", x"0f21", x"0f21", x"0f21", x"0f21", x"0f21", x"0f21", x"0f21", x"0f21", x"0f21", x"0f21", x"0f21", x"0f21", x"0f21", x"0f22", x"0f22", x"0f22", x"0f22", x"0f22", x"0f22", x"0f22", x"0f22", x"0f22", x"0f22", x"0f22", x"0f22", x"0f22", x"0f22", x"0f22", x"0f22", x"0f22", x"0f22", x"0f22", x"0f22", x"0f23", x"0f23", x"0f23", x"0f23", x"0f23", x"0f23", x"0f23", x"0f23", x"0f23", x"0f23", x"0f23", x"0f23", x"0f23", x"0f23", x"0f23", x"0f23", x"0f23", x"0f23", x"0f23", x"0f24", x"0f24", x"0f24", x"0f24", x"0f24", x"0f24", x"0f24", x"0f24", x"0f24", x"0f24", x"0f24", x"0f24", x"0f24", x"0f24", x"0f24", x"0f24", x"0f24", x"0f24", x"0f24", x"0f24", x"0f25", x"0f25", x"0f25", x"0f25", x"0f25", x"0f25", x"0f25", x"0f25", x"0f25", x"0f25", x"0f25", x"0f25", x"0f25", x"0f25", x"0f25", x"0f25", x"0f25", x"0f25", x"0f25", x"0f25", x"0f26", x"0f26", x"0f26", x"0f26", x"0f26", x"0f26", x"0f26", x"0f26", x"0f26", x"0f26", x"0f26", x"0f26", x"0f26", x"0f26", x"0f26", x"0f26", x"0f26", x"0f26", x"0f26", x"0f26", x"0f27", x"0f27", x"0f27", x"0f27", x"0f27", x"0f27", x"0f27", x"0f27", x"0f27", x"0f27", x"0f27", x"0f27", x"0f27", x"0f27", x"0f27", x"0f27", x"0f27", x"0f27", x"0f27", x"0f27", x"0f28", x"0f28", x"0f28", x"0f28", x"0f28", x"0f28", x"0f28", x"0f28", x"0f28", x"0f28", x"0f28", x"0f28", x"0f28", x"0f28", x"0f28", x"0f28", x"0f28", x"0f28", x"0f28", x"0f28", x"0f29", x"0f29", x"0f29", x"0f29", x"0f29", x"0f29", x"0f29", x"0f29", x"0f29", x"0f29", x"0f29", x"0f29", x"0f29", x"0f29", x"0f29", x"0f29", x"0f29", x"0f29", x"0f29", x"0f29", x"0f2a", x"0f2a", x"0f2a", x"0f2a", x"0f2a", x"0f2a", x"0f2a", x"0f2a", x"0f2a", x"0f2a", x"0f2a", x"0f2a", x"0f2a", x"0f2a", x"0f2a", x"0f2a", x"0f2a", x"0f2a", x"0f2a", x"0f2a", x"0f2a", x"0f2b", x"0f2b", x"0f2b", x"0f2b", x"0f2b", x"0f2b", x"0f2b", x"0f2b", x"0f2b", x"0f2b", x"0f2b", x"0f2b", x"0f2b", x"0f2b", x"0f2b", x"0f2b", x"0f2b", x"0f2b", x"0f2b", x"0f2b", x"0f2c", x"0f2c", x"0f2c", x"0f2c", x"0f2c", x"0f2c", x"0f2c", x"0f2c", x"0f2c", x"0f2c", x"0f2c", x"0f2c", x"0f2c", x"0f2c", x"0f2c", x"0f2c", x"0f2c", x"0f2c", x"0f2c", x"0f2c", x"0f2c", x"0f2d", x"0f2d", x"0f2d", x"0f2d", x"0f2d", x"0f2d", x"0f2d", x"0f2d", x"0f2d", x"0f2d", x"0f2d", x"0f2d", x"0f2d", x"0f2d", x"0f2d", x"0f2d", x"0f2d", x"0f2d", x"0f2d", x"0f2d", x"0f2e", x"0f2e", x"0f2e", x"0f2e", x"0f2e", x"0f2e", x"0f2e", x"0f2e", x"0f2e", x"0f2e", x"0f2e", x"0f2e", x"0f2e", x"0f2e", x"0f2e", x"0f2e", x"0f2e", x"0f2e", x"0f2e", x"0f2e", x"0f2e", x"0f2f", x"0f2f", x"0f2f", x"0f2f", x"0f2f", x"0f2f", x"0f2f", x"0f2f", x"0f2f", x"0f2f", x"0f2f", x"0f2f", x"0f2f", x"0f2f", x"0f2f", x"0f2f", x"0f2f", x"0f2f", x"0f2f", x"0f2f", x"0f2f", x"0f30", x"0f30", x"0f30", x"0f30", x"0f30", x"0f30", x"0f30", x"0f30", x"0f30", x"0f30", x"0f30", x"0f30", x"0f30", x"0f30", x"0f30", x"0f30", x"0f30", x"0f30", x"0f30", x"0f30", x"0f30", x"0f31", x"0f31", x"0f31", x"0f31", x"0f31", x"0f31", x"0f31", x"0f31", x"0f31", x"0f31", x"0f31", x"0f31", x"0f31", x"0f31", x"0f31", x"0f31", x"0f31", x"0f31", x"0f31", x"0f31", x"0f31", x"0f32", x"0f32", x"0f32", x"0f32", x"0f32", x"0f32", x"0f32", x"0f32", x"0f32", x"0f32", x"0f32", x"0f32", x"0f32", x"0f32", x"0f32", x"0f32", x"0f32", x"0f32", x"0f32", x"0f32", x"0f32", x"0f33", x"0f33", x"0f33", x"0f33", x"0f33", x"0f33", x"0f33", x"0f33", x"0f33", x"0f33", x"0f33", x"0f33", x"0f33", x"0f33", x"0f33", x"0f33", x"0f33", x"0f33", x"0f33", x"0f33", x"0f33", x"0f34", x"0f34", x"0f34", x"0f34", x"0f34", x"0f34", x"0f34", x"0f34", x"0f34", x"0f34", x"0f34", x"0f34", x"0f34", x"0f34", x"0f34", x"0f34", x"0f34", x"0f34", x"0f34", x"0f34", x"0f34", x"0f35", x"0f35", x"0f35", x"0f35", x"0f35", x"0f35", x"0f35", x"0f35", x"0f35", x"0f35", x"0f35", x"0f35", x"0f35", x"0f35", x"0f35", x"0f35", x"0f35", x"0f35", x"0f35", x"0f35", x"0f35", x"0f35", x"0f36", x"0f36", x"0f36", x"0f36", x"0f36", x"0f36", x"0f36", x"0f36", x"0f36", x"0f36", x"0f36", x"0f36", x"0f36", x"0f36", x"0f36", x"0f36", x"0f36", x"0f36", x"0f36", x"0f36", x"0f36", x"0f37", x"0f37", x"0f37", x"0f37", x"0f37", x"0f37", x"0f37", x"0f37", x"0f37", x"0f37", x"0f37", x"0f37", x"0f37", x"0f37", x"0f37", x"0f37", x"0f37", x"0f37", x"0f37", x"0f37", x"0f37", x"0f37", x"0f38", x"0f38", x"0f38", x"0f38", x"0f38", x"0f38", x"0f38", x"0f38", x"0f38", x"0f38", x"0f38", x"0f38", x"0f38", x"0f38", x"0f38", x"0f38", x"0f38", x"0f38", x"0f38", x"0f38", x"0f38", x"0f39", x"0f39", x"0f39", x"0f39", x"0f39", x"0f39", x"0f39", x"0f39", x"0f39", x"0f39", x"0f39", x"0f39", x"0f39", x"0f39", x"0f39", x"0f39", x"0f39", x"0f39", x"0f39", x"0f39", x"0f39", x"0f39", x"0f3a", x"0f3a", x"0f3a", x"0f3a", x"0f3a", x"0f3a", x"0f3a", x"0f3a", x"0f3a", x"0f3a", x"0f3a", x"0f3a", x"0f3a", x"0f3a", x"0f3a", x"0f3a", x"0f3a", x"0f3a", x"0f3a", x"0f3a", x"0f3a", x"0f3a", x"0f3b", x"0f3b", x"0f3b", x"0f3b", x"0f3b", x"0f3b", x"0f3b", x"0f3b", x"0f3b", x"0f3b", x"0f3b", x"0f3b", x"0f3b", x"0f3b", x"0f3b", x"0f3b", x"0f3b", x"0f3b", x"0f3b", x"0f3b", x"0f3b", x"0f3b", x"0f3c", x"0f3c", x"0f3c", x"0f3c", x"0f3c", x"0f3c", x"0f3c", x"0f3c", x"0f3c", x"0f3c", x"0f3c", x"0f3c", x"0f3c", x"0f3c", x"0f3c", x"0f3c", x"0f3c", x"0f3c", x"0f3c", x"0f3c", x"0f3c", x"0f3c", x"0f3d", x"0f3d", x"0f3d", x"0f3d", x"0f3d", x"0f3d", x"0f3d", x"0f3d", x"0f3d", x"0f3d", x"0f3d", x"0f3d", x"0f3d", x"0f3d", x"0f3d", x"0f3d", x"0f3d", x"0f3d", x"0f3d", x"0f3d", x"0f3d", x"0f3d", x"0f3e", x"0f3e", x"0f3e", x"0f3e", x"0f3e", x"0f3e", x"0f3e", x"0f3e", x"0f3e", x"0f3e", x"0f3e", x"0f3e", x"0f3e", x"0f3e", x"0f3e", x"0f3e", x"0f3e", x"0f3e", x"0f3e", x"0f3e", x"0f3e", x"0f3e", x"0f3e", x"0f3f", x"0f3f", x"0f3f", x"0f3f", x"0f3f", x"0f3f", x"0f3f", x"0f3f", x"0f3f", x"0f3f", x"0f3f", x"0f3f", x"0f3f", x"0f3f", x"0f3f", x"0f3f", x"0f3f", x"0f3f", x"0f3f", x"0f3f", x"0f3f", x"0f3f", x"0f40", x"0f40", x"0f40", x"0f40", x"0f40", x"0f40", x"0f40", x"0f40", x"0f40", x"0f40", x"0f40", x"0f40", x"0f40", x"0f40", x"0f40", x"0f40", x"0f40", x"0f40", x"0f40", x"0f40", x"0f40", x"0f40", x"0f40", x"0f41", x"0f41", x"0f41", x"0f41", x"0f41", x"0f41", x"0f41", x"0f41", x"0f41", x"0f41", x"0f41", x"0f41", x"0f41", x"0f41", x"0f41", x"0f41", x"0f41", x"0f41", x"0f41", x"0f41", x"0f41", x"0f41", x"0f42", x"0f42", x"0f42", x"0f42", x"0f42", x"0f42", x"0f42", x"0f42", x"0f42", x"0f42", x"0f42", x"0f42", x"0f42", x"0f42", x"0f42", x"0f42", x"0f42", x"0f42", x"0f42", x"0f42", x"0f42", x"0f42", x"0f42", x"0f43", x"0f43", x"0f43", x"0f43", x"0f43", x"0f43", x"0f43", x"0f43", x"0f43", x"0f43", x"0f43", x"0f43", x"0f43", x"0f43", x"0f43", x"0f43", x"0f43", x"0f43", x"0f43", x"0f43", x"0f43", x"0f43", x"0f43", x"0f44", x"0f44", x"0f44", x"0f44", x"0f44", x"0f44", x"0f44", x"0f44", x"0f44", x"0f44", x"0f44", x"0f44", x"0f44", x"0f44", x"0f44", x"0f44", x"0f44", x"0f44", x"0f44", x"0f44", x"0f44", x"0f44", x"0f44", x"0f45", x"0f45", x"0f45", x"0f45", x"0f45", x"0f45", x"0f45", x"0f45", x"0f45", x"0f45", x"0f45", x"0f45", x"0f45", x"0f45", x"0f45", x"0f45", x"0f45", x"0f45", x"0f45", x"0f45", x"0f45", x"0f45", x"0f45", x"0f46", x"0f46", x"0f46", x"0f46", x"0f46", x"0f46", x"0f46", x"0f46", x"0f46", x"0f46", x"0f46", x"0f46", x"0f46", x"0f46", x"0f46", x"0f46", x"0f46", x"0f46", x"0f46", x"0f46", x"0f46", x"0f46", x"0f46", x"0f47", x"0f47", x"0f47", x"0f47", x"0f47", x"0f47", x"0f47", x"0f47", x"0f47", x"0f47", x"0f47", x"0f47", x"0f47", x"0f47", x"0f47", x"0f47", x"0f47", x"0f47", x"0f47", x"0f47", x"0f47", x"0f47", x"0f47", x"0f47", x"0f48", x"0f48", x"0f48", x"0f48", x"0f48", x"0f48", x"0f48", x"0f48", x"0f48", x"0f48", x"0f48", x"0f48", x"0f48", x"0f48", x"0f48", x"0f48", x"0f48", x"0f48", x"0f48", x"0f48", x"0f48", x"0f48", x"0f48", x"0f49", x"0f49", x"0f49", x"0f49", x"0f49", x"0f49", x"0f49", x"0f49", x"0f49", x"0f49", x"0f49", x"0f49", x"0f49", x"0f49", x"0f49", x"0f49", x"0f49", x"0f49", x"0f49", x"0f49", x"0f49", x"0f49", x"0f49", x"0f49", x"0f4a", x"0f4a", x"0f4a", x"0f4a", x"0f4a", x"0f4a", x"0f4a", x"0f4a", x"0f4a", x"0f4a", x"0f4a", x"0f4a", x"0f4a", x"0f4a", x"0f4a", x"0f4a", x"0f4a", x"0f4a", x"0f4a", x"0f4a", x"0f4a", x"0f4a", x"0f4a", x"0f4a", x"0f4b", x"0f4b", x"0f4b", x"0f4b", x"0f4b", x"0f4b", x"0f4b", x"0f4b", x"0f4b", x"0f4b", x"0f4b", x"0f4b", x"0f4b", x"0f4b", x"0f4b", x"0f4b", x"0f4b", x"0f4b", x"0f4b", x"0f4b", x"0f4b", x"0f4b", x"0f4b", x"0f4c", x"0f4c", x"0f4c", x"0f4c", x"0f4c", x"0f4c", x"0f4c", x"0f4c", x"0f4c", x"0f4c", x"0f4c", x"0f4c", x"0f4c", x"0f4c", x"0f4c", x"0f4c", x"0f4c", x"0f4c", x"0f4c", x"0f4c", x"0f4c", x"0f4c", x"0f4c", x"0f4c", x"0f4d", x"0f4d", x"0f4d", x"0f4d", x"0f4d", x"0f4d", x"0f4d", x"0f4d", x"0f4d", x"0f4d", x"0f4d", x"0f4d", x"0f4d", x"0f4d", x"0f4d", x"0f4d", x"0f4d", x"0f4d", x"0f4d", x"0f4d", x"0f4d", x"0f4d", x"0f4d", x"0f4d", x"0f4d", x"0f4e", x"0f4e", x"0f4e", x"0f4e", x"0f4e", x"0f4e", x"0f4e", x"0f4e", x"0f4e", x"0f4e", x"0f4e", x"0f4e", x"0f4e", x"0f4e", x"0f4e", x"0f4e", x"0f4e", x"0f4e", x"0f4e", x"0f4e", x"0f4e", x"0f4e", x"0f4e", x"0f4e", x"0f4f", x"0f4f", x"0f4f", x"0f4f", x"0f4f", x"0f4f", x"0f4f", x"0f4f", x"0f4f", x"0f4f", x"0f4f", x"0f4f", x"0f4f", x"0f4f", x"0f4f", x"0f4f", x"0f4f", x"0f4f", x"0f4f", x"0f4f", x"0f4f", x"0f4f", x"0f4f", x"0f4f", x"0f50", x"0f50", x"0f50", x"0f50", x"0f50", x"0f50", x"0f50", x"0f50", x"0f50", x"0f50", x"0f50", x"0f50", x"0f50", x"0f50", x"0f50", x"0f50", x"0f50", x"0f50", x"0f50", x"0f50", x"0f50", x"0f50", x"0f50", x"0f50", x"0f50", x"0f51", x"0f51", x"0f51", x"0f51", x"0f51", x"0f51", x"0f51", x"0f51", x"0f51", x"0f51", x"0f51", x"0f51", x"0f51", x"0f51", x"0f51", x"0f51", x"0f51", x"0f51", x"0f51", x"0f51", x"0f51", x"0f51", x"0f51", x"0f51", x"0f52", x"0f52", x"0f52", x"0f52", x"0f52", x"0f52", x"0f52", x"0f52", x"0f52", x"0f52", x"0f52", x"0f52", x"0f52", x"0f52", x"0f52", x"0f52", x"0f52", x"0f52", x"0f52", x"0f52", x"0f52", x"0f52", x"0f52", x"0f52", x"0f52", x"0f53", x"0f53", x"0f53", x"0f53", x"0f53", x"0f53", x"0f53", x"0f53", x"0f53", x"0f53", x"0f53", x"0f53", x"0f53", x"0f53", x"0f53", x"0f53", x"0f53", x"0f53", x"0f53", x"0f53", x"0f53", x"0f53", x"0f53", x"0f53", x"0f53", x"0f54", x"0f54", x"0f54", x"0f54", x"0f54", x"0f54", x"0f54", x"0f54", x"0f54", x"0f54", x"0f54", x"0f54", x"0f54", x"0f54", x"0f54", x"0f54", x"0f54", x"0f54", x"0f54", x"0f54", x"0f54", x"0f54", x"0f54", x"0f54", x"0f54", x"0f55", x"0f55", x"0f55", x"0f55", x"0f55", x"0f55", x"0f55", x"0f55", x"0f55", x"0f55", x"0f55", x"0f55", x"0f55", x"0f55", x"0f55", x"0f55", x"0f55", x"0f55", x"0f55", x"0f55", x"0f55", x"0f55", x"0f55", x"0f55", x"0f55", x"0f56", x"0f56", x"0f56", x"0f56", x"0f56", x"0f56", x"0f56", x"0f56", x"0f56", x"0f56", x"0f56", x"0f56", x"0f56", x"0f56", x"0f56", x"0f56", x"0f56", x"0f56", x"0f56", x"0f56", x"0f56", x"0f56", x"0f56", x"0f56", x"0f56", x"0f56", x"0f57", x"0f57", x"0f57", x"0f57", x"0f57", x"0f57", x"0f57", x"0f57", x"0f57", x"0f57", x"0f57", x"0f57", x"0f57", x"0f57", x"0f57", x"0f57", x"0f57", x"0f57", x"0f57", x"0f57", x"0f57", x"0f57", x"0f57", x"0f57", x"0f57", x"0f58", x"0f58", x"0f58", x"0f58", x"0f58", x"0f58", x"0f58", x"0f58", x"0f58", x"0f58", x"0f58", x"0f58", x"0f58", x"0f58", x"0f58", x"0f58", x"0f58", x"0f58", x"0f58", x"0f58", x"0f58", x"0f58", x"0f58", x"0f58", x"0f58", x"0f58", x"0f59", x"0f59", x"0f59", x"0f59", x"0f59", x"0f59", x"0f59", x"0f59", x"0f59", x"0f59", x"0f59", x"0f59", x"0f59", x"0f59", x"0f59", x"0f59", x"0f59", x"0f59", x"0f59", x"0f59", x"0f59", x"0f59", x"0f59", x"0f59", x"0f59", x"0f59", x"0f5a", x"0f5a", x"0f5a", x"0f5a", x"0f5a", x"0f5a", x"0f5a", x"0f5a", x"0f5a", x"0f5a", x"0f5a", x"0f5a", x"0f5a", x"0f5a", x"0f5a", x"0f5a", x"0f5a", x"0f5a", x"0f5a", x"0f5a", x"0f5a", x"0f5a", x"0f5a", x"0f5a", x"0f5a", x"0f5a", x"0f5b", x"0f5b", x"0f5b", x"0f5b", x"0f5b", x"0f5b", x"0f5b", x"0f5b", x"0f5b", x"0f5b", x"0f5b", x"0f5b", x"0f5b", x"0f5b", x"0f5b", x"0f5b", x"0f5b", x"0f5b", x"0f5b", x"0f5b", x"0f5b", x"0f5b", x"0f5b", x"0f5b", x"0f5b", x"0f5b", x"0f5c", x"0f5c", x"0f5c", x"0f5c", x"0f5c", x"0f5c", x"0f5c", x"0f5c", x"0f5c", x"0f5c", x"0f5c", x"0f5c", x"0f5c", x"0f5c", x"0f5c", x"0f5c", x"0f5c", x"0f5c", x"0f5c", x"0f5c", x"0f5c", x"0f5c", x"0f5c", x"0f5c", x"0f5c", x"0f5c", x"0f5d", x"0f5d", x"0f5d", x"0f5d", x"0f5d", x"0f5d", x"0f5d", x"0f5d", x"0f5d", x"0f5d", x"0f5d", x"0f5d", x"0f5d", x"0f5d", x"0f5d", x"0f5d", x"0f5d", x"0f5d", x"0f5d", x"0f5d", x"0f5d", x"0f5d", x"0f5d", x"0f5d", x"0f5d", x"0f5d", x"0f5e", x"0f5e", x"0f5e", x"0f5e", x"0f5e", x"0f5e", x"0f5e", x"0f5e", x"0f5e", x"0f5e", x"0f5e", x"0f5e", x"0f5e", x"0f5e", x"0f5e", x"0f5e", x"0f5e", x"0f5e", x"0f5e", x"0f5e", x"0f5e", x"0f5e", x"0f5e", x"0f5e", x"0f5e", x"0f5e", x"0f5e", x"0f5f", x"0f5f", x"0f5f", x"0f5f", x"0f5f", x"0f5f", x"0f5f", x"0f5f", x"0f5f", x"0f5f", x"0f5f", x"0f5f", x"0f5f", x"0f5f", x"0f5f", x"0f5f", x"0f5f", x"0f5f", x"0f5f", x"0f5f", x"0f5f", x"0f5f", x"0f5f", x"0f5f", x"0f5f", x"0f5f", x"0f5f", x"0f60", x"0f60", x"0f60", x"0f60", x"0f60", x"0f60", x"0f60", x"0f60", x"0f60", x"0f60", x"0f60", x"0f60", x"0f60", x"0f60", x"0f60", x"0f60", x"0f60", x"0f60", x"0f60", x"0f60", x"0f60", x"0f60", x"0f60", x"0f60", x"0f60", x"0f60", x"0f60", x"0f61", x"0f61", x"0f61", x"0f61", x"0f61", x"0f61", x"0f61", x"0f61", x"0f61", x"0f61", x"0f61", x"0f61", x"0f61", x"0f61", x"0f61", x"0f61", x"0f61", x"0f61", x"0f61", x"0f61", x"0f61", x"0f61", x"0f61", x"0f61", x"0f61", x"0f61", x"0f61", x"0f62", x"0f62", x"0f62", x"0f62", x"0f62", x"0f62", x"0f62", x"0f62", x"0f62", x"0f62", x"0f62", x"0f62", x"0f62", x"0f62", x"0f62", x"0f62", x"0f62", x"0f62", x"0f62", x"0f62", x"0f62", x"0f62", x"0f62", x"0f62", x"0f62", x"0f62", x"0f62", x"0f63", x"0f63", x"0f63", x"0f63", x"0f63", x"0f63", x"0f63", x"0f63", x"0f63", x"0f63", x"0f63", x"0f63", x"0f63", x"0f63", x"0f63", x"0f63", x"0f63", x"0f63", x"0f63", x"0f63", x"0f63", x"0f63", x"0f63", x"0f63", x"0f63", x"0f63", x"0f63", x"0f64", x"0f64", x"0f64", x"0f64", x"0f64", x"0f64", x"0f64", x"0f64", x"0f64", x"0f64", x"0f64", x"0f64", x"0f64", x"0f64", x"0f64", x"0f64", x"0f64", x"0f64", x"0f64", x"0f64", x"0f64", x"0f64", x"0f64", x"0f64", x"0f64", x"0f64", x"0f64", x"0f64", x"0f65", x"0f65", x"0f65", x"0f65", x"0f65", x"0f65", x"0f65", x"0f65", x"0f65", x"0f65", x"0f65", x"0f65", x"0f65", x"0f65", x"0f65", x"0f65", x"0f65", x"0f65", x"0f65", x"0f65", x"0f65", x"0f65", x"0f65", x"0f65", x"0f65", x"0f65", x"0f65", x"0f66", x"0f66", x"0f66", x"0f66", x"0f66", x"0f66", x"0f66", x"0f66", x"0f66", x"0f66", x"0f66", x"0f66", x"0f66", x"0f66", x"0f66", x"0f66", x"0f66", x"0f66", x"0f66", x"0f66", x"0f66", x"0f66", x"0f66", x"0f66", x"0f66", x"0f66", x"0f66", x"0f66", x"0f67", x"0f67", x"0f67", x"0f67", x"0f67", x"0f67", x"0f67", x"0f67", x"0f67", x"0f67", x"0f67", x"0f67", x"0f67", x"0f67", x"0f67", x"0f67", x"0f67", x"0f67", x"0f67", x"0f67", x"0f67", x"0f67", x"0f67", x"0f67", x"0f67", x"0f67", x"0f67", x"0f67", x"0f68", x"0f68", x"0f68", x"0f68", x"0f68", x"0f68", x"0f68", x"0f68", x"0f68", x"0f68", x"0f68", x"0f68", x"0f68", x"0f68", x"0f68", x"0f68", x"0f68", x"0f68", x"0f68", x"0f68", x"0f68", x"0f68", x"0f68", x"0f68", x"0f68", x"0f68", x"0f68", x"0f68", x"0f68", x"0f69", x"0f69", x"0f69", x"0f69", x"0f69", x"0f69", x"0f69", x"0f69", x"0f69", x"0f69", x"0f69", x"0f69", x"0f69", x"0f69", x"0f69", x"0f69", x"0f69", x"0f69", x"0f69", x"0f69", x"0f69", x"0f69", x"0f69", x"0f69", x"0f69", x"0f69", x"0f69", x"0f69", x"0f6a", x"0f6a", x"0f6a", x"0f6a", x"0f6a", x"0f6a", x"0f6a", x"0f6a", x"0f6a", x"0f6a", x"0f6a", x"0f6a", x"0f6a", x"0f6a", x"0f6a", x"0f6a", x"0f6a", x"0f6a", x"0f6a", x"0f6a", x"0f6a", x"0f6a", x"0f6a", x"0f6a", x"0f6a", x"0f6a", x"0f6a", x"0f6a", x"0f6a", x"0f6b", x"0f6b", x"0f6b", x"0f6b", x"0f6b", x"0f6b", x"0f6b", x"0f6b", x"0f6b", x"0f6b", x"0f6b", x"0f6b", x"0f6b", x"0f6b", x"0f6b", x"0f6b", x"0f6b", x"0f6b", x"0f6b", x"0f6b", x"0f6b", x"0f6b", x"0f6b", x"0f6b", x"0f6b", x"0f6b", x"0f6b", x"0f6b", x"0f6b", x"0f6c", x"0f6c", x"0f6c", x"0f6c", x"0f6c", x"0f6c", x"0f6c", x"0f6c", x"0f6c", x"0f6c", x"0f6c", x"0f6c", x"0f6c", x"0f6c", x"0f6c", x"0f6c", x"0f6c", x"0f6c", x"0f6c", x"0f6c", x"0f6c", x"0f6c", x"0f6c", x"0f6c", x"0f6c", x"0f6c", x"0f6c", x"0f6c", x"0f6c", x"0f6d", x"0f6d", x"0f6d", x"0f6d", x"0f6d", x"0f6d", x"0f6d", x"0f6d", x"0f6d", x"0f6d", x"0f6d", x"0f6d", x"0f6d", x"0f6d", x"0f6d", x"0f6d", x"0f6d", x"0f6d", x"0f6d", x"0f6d", x"0f6d", x"0f6d", x"0f6d", x"0f6d", x"0f6d", x"0f6d", x"0f6d", x"0f6d", x"0f6d", x"0f6e", x"0f6e", x"0f6e", x"0f6e", x"0f6e", x"0f6e", x"0f6e", x"0f6e", x"0f6e", x"0f6e", x"0f6e", x"0f6e", x"0f6e", x"0f6e", x"0f6e", x"0f6e", x"0f6e", x"0f6e", x"0f6e", x"0f6e", x"0f6e", x"0f6e", x"0f6e", x"0f6e", x"0f6e", x"0f6e", x"0f6e", x"0f6e", x"0f6e", x"0f6f", x"0f6f", x"0f6f", x"0f6f", x"0f6f", x"0f6f", x"0f6f", x"0f6f", x"0f6f", x"0f6f", x"0f6f", x"0f6f", x"0f6f", x"0f6f", x"0f6f", x"0f6f", x"0f6f", x"0f6f", x"0f6f", x"0f6f", x"0f6f", x"0f6f", x"0f6f", x"0f6f", x"0f6f", x"0f6f", x"0f6f", x"0f6f", x"0f6f", x"0f6f", x"0f70", x"0f70", x"0f70", x"0f70", x"0f70", x"0f70", x"0f70", x"0f70", x"0f70", x"0f70", x"0f70", x"0f70", x"0f70", x"0f70", x"0f70", x"0f70", x"0f70", x"0f70", x"0f70", x"0f70", x"0f70", x"0f70", x"0f70", x"0f70", x"0f70", x"0f70", x"0f70", x"0f70", x"0f70", x"0f71", x"0f71", x"0f71", x"0f71", x"0f71", x"0f71", x"0f71", x"0f71", x"0f71", x"0f71", x"0f71", x"0f71", x"0f71", x"0f71", x"0f71", x"0f71", x"0f71", x"0f71", x"0f71", x"0f71", x"0f71", x"0f71", x"0f71", x"0f71", x"0f71", x"0f71", x"0f71", x"0f71", x"0f71", x"0f71", x"0f72", x"0f72", x"0f72", x"0f72", x"0f72", x"0f72", x"0f72", x"0f72", x"0f72", x"0f72", x"0f72", x"0f72", x"0f72", x"0f72", x"0f72", x"0f72", x"0f72", x"0f72", x"0f72", x"0f72", x"0f72", x"0f72", x"0f72", x"0f72", x"0f72", x"0f72", x"0f72", x"0f72", x"0f72", x"0f72", x"0f72", x"0f73", x"0f73", x"0f73", x"0f73", x"0f73", x"0f73", x"0f73", x"0f73", x"0f73", x"0f73", x"0f73", x"0f73", x"0f73", x"0f73", x"0f73", x"0f73", x"0f73", x"0f73", x"0f73", x"0f73", x"0f73", x"0f73", x"0f73", x"0f73", x"0f73", x"0f73", x"0f73", x"0f73", x"0f73", x"0f73", x"0f74", x"0f74", x"0f74", x"0f74", x"0f74", x"0f74", x"0f74", x"0f74", x"0f74", x"0f74", x"0f74", x"0f74", x"0f74", x"0f74", x"0f74", x"0f74", x"0f74", x"0f74", x"0f74", x"0f74", x"0f74", x"0f74", x"0f74", x"0f74", x"0f74", x"0f74", x"0f74", x"0f74", x"0f74", x"0f74", x"0f74", x"0f75", x"0f75", x"0f75", x"0f75", x"0f75", x"0f75", x"0f75", x"0f75", x"0f75", x"0f75", x"0f75", x"0f75", x"0f75", x"0f75", x"0f75", x"0f75", x"0f75", x"0f75", x"0f75", x"0f75", x"0f75", x"0f75", x"0f75", x"0f75", x"0f75", x"0f75", x"0f75", x"0f75", x"0f75", x"0f75", x"0f76", x"0f76", x"0f76", x"0f76", x"0f76", x"0f76", x"0f76", x"0f76", x"0f76", x"0f76", x"0f76", x"0f76", x"0f76", x"0f76", x"0f76", x"0f76", x"0f76", x"0f76", x"0f76", x"0f76", x"0f76", x"0f76", x"0f76", x"0f76", x"0f76", x"0f76", x"0f76", x"0f76", x"0f76", x"0f76", x"0f76", x"0f77", x"0f77", x"0f77", x"0f77", x"0f77", x"0f77", x"0f77", x"0f77", x"0f77", x"0f77", x"0f77", x"0f77", x"0f77", x"0f77", x"0f77", x"0f77", x"0f77", x"0f77", x"0f77", x"0f77", x"0f77", x"0f77", x"0f77", x"0f77", x"0f77", x"0f77", x"0f77", x"0f77", x"0f77", x"0f77", x"0f77", x"0f77", x"0f78", x"0f78", x"0f78", x"0f78", x"0f78", x"0f78", x"0f78", x"0f78", x"0f78", x"0f78", x"0f78", x"0f78", x"0f78", x"0f78", x"0f78", x"0f78", x"0f78", x"0f78", x"0f78", x"0f78", x"0f78", x"0f78", x"0f78", x"0f78", x"0f78", x"0f78", x"0f78", x"0f78", x"0f78", x"0f78", x"0f78", x"0f79", x"0f79", x"0f79", x"0f79", x"0f79", x"0f79", x"0f79", x"0f79", x"0f79", x"0f79", x"0f79", x"0f79", x"0f79", x"0f79", x"0f79", x"0f79", x"0f79", x"0f79", x"0f79", x"0f79", x"0f79", x"0f79", x"0f79", x"0f79", x"0f79", x"0f79", x"0f79", x"0f79", x"0f79", x"0f79", x"0f79", x"0f79", x"0f7a", x"0f7a", x"0f7a", x"0f7a", x"0f7a", x"0f7a", x"0f7a", x"0f7a", x"0f7a", x"0f7a", x"0f7a", x"0f7a", x"0f7a", x"0f7a", x"0f7a", x"0f7a", x"0f7a", x"0f7a", x"0f7a", x"0f7a", x"0f7a", x"0f7a", x"0f7a", x"0f7a", x"0f7a", x"0f7a", x"0f7a", x"0f7a", x"0f7a", x"0f7a", x"0f7a", x"0f7a", x"0f7b", x"0f7b", x"0f7b", x"0f7b", x"0f7b", x"0f7b", x"0f7b", x"0f7b", x"0f7b", x"0f7b", x"0f7b", x"0f7b", x"0f7b", x"0f7b", x"0f7b", x"0f7b", x"0f7b", x"0f7b", x"0f7b", x"0f7b", x"0f7b", x"0f7b", x"0f7b", x"0f7b", x"0f7b", x"0f7b", x"0f7b", x"0f7b", x"0f7b", x"0f7b", x"0f7b", x"0f7b", x"0f7c", x"0f7c", x"0f7c", x"0f7c", x"0f7c", x"0f7c", x"0f7c", x"0f7c", x"0f7c", x"0f7c", x"0f7c", x"0f7c", x"0f7c", x"0f7c", x"0f7c", x"0f7c", x"0f7c", x"0f7c", x"0f7c", x"0f7c", x"0f7c", x"0f7c", x"0f7c", x"0f7c", x"0f7c", x"0f7c", x"0f7c", x"0f7c", x"0f7c", x"0f7c", x"0f7c", x"0f7c", x"0f7c", x"0f7d", x"0f7d", x"0f7d", x"0f7d", x"0f7d", x"0f7d", x"0f7d", x"0f7d", x"0f7d", x"0f7d", x"0f7d", x"0f7d", x"0f7d", x"0f7d", x"0f7d", x"0f7d", x"0f7d", x"0f7d", x"0f7d", x"0f7d", x"0f7d", x"0f7d", x"0f7d", x"0f7d", x"0f7d", x"0f7d", x"0f7d", x"0f7d", x"0f7d", x"0f7d", x"0f7d", x"0f7d", x"0f7e", x"0f7e", x"0f7e", x"0f7e", x"0f7e", x"0f7e", x"0f7e", x"0f7e", x"0f7e", x"0f7e", x"0f7e", x"0f7e", x"0f7e", x"0f7e", x"0f7e", x"0f7e", x"0f7e", x"0f7e", x"0f7e", x"0f7e", x"0f7e", x"0f7e", x"0f7e", x"0f7e", x"0f7e", x"0f7e", x"0f7e", x"0f7e", x"0f7e", x"0f7e", x"0f7e", x"0f7e", x"0f7e", x"0f7f", x"0f7f", x"0f7f", x"0f7f", x"0f7f", x"0f7f", x"0f7f", x"0f7f", x"0f7f", x"0f7f", x"0f7f", x"0f7f", x"0f7f", x"0f7f", x"0f7f", x"0f7f", x"0f7f", x"0f7f", x"0f7f", x"0f7f", x"0f7f", x"0f7f", x"0f7f", x"0f7f", x"0f7f", x"0f7f", x"0f7f", x"0f7f", x"0f7f", x"0f7f", x"0f7f", x"0f7f", x"0f7f", x"0f80", x"0f80", x"0f80", x"0f80", x"0f80", x"0f80", x"0f80", x"0f80", x"0f80", x"0f80", x"0f80", x"0f80", x"0f80", x"0f80", x"0f80", x"0f80", x"0f80", x"0f80", x"0f80", x"0f80", x"0f80", x"0f80", x"0f80", x"0f80", x"0f80", x"0f80", x"0f80", x"0f80", x"0f80", x"0f80", x"0f80", x"0f80", x"0f80", x"0f80", x"0f81", x"0f81", x"0f81", x"0f81", x"0f81", x"0f81", x"0f81", x"0f81", x"0f81", x"0f81", x"0f81", x"0f81", x"0f81", x"0f81", x"0f81", x"0f81", x"0f81", x"0f81", x"0f81", x"0f81", x"0f81", x"0f81", x"0f81", x"0f81", x"0f81", x"0f81", x"0f81", x"0f81", x"0f81", x"0f81", x"0f81", x"0f81", x"0f81", x"0f82", x"0f82", x"0f82", x"0f82", x"0f82", x"0f82", x"0f82", x"0f82", x"0f82", x"0f82", x"0f82", x"0f82", x"0f82", x"0f82", x"0f82", x"0f82", x"0f82", x"0f82", x"0f82", x"0f82", x"0f82", x"0f82", x"0f82", x"0f82", x"0f82", x"0f82", x"0f82", x"0f82", x"0f82", x"0f82", x"0f82", x"0f82", x"0f82", x"0f82", x"0f83", x"0f83", x"0f83", x"0f83", x"0f83", x"0f83", x"0f83", x"0f83", x"0f83", x"0f83", x"0f83", x"0f83", x"0f83", x"0f83", x"0f83", x"0f83", x"0f83", x"0f83", x"0f83", x"0f83", x"0f83", x"0f83", x"0f83", x"0f83", x"0f83", x"0f83", x"0f83", x"0f83", x"0f83", x"0f83", x"0f83", x"0f83", x"0f83", x"0f83", x"0f84", x"0f84", x"0f84", x"0f84", x"0f84", x"0f84", x"0f84", x"0f84", x"0f84", x"0f84", x"0f84", x"0f84", x"0f84", x"0f84", x"0f84", x"0f84", x"0f84", x"0f84", x"0f84", x"0f84", x"0f84", x"0f84", x"0f84", x"0f84", x"0f84", x"0f84", x"0f84", x"0f84", x"0f84", x"0f84", x"0f84", x"0f84", x"0f84", x"0f84", x"0f84", x"0f85", x"0f85", x"0f85", x"0f85", x"0f85", x"0f85", x"0f85", x"0f85", x"0f85", x"0f85", x"0f85", x"0f85", x"0f85", x"0f85", x"0f85", x"0f85", x"0f85", x"0f85", x"0f85", x"0f85", x"0f85", x"0f85", x"0f85", x"0f85", x"0f85", x"0f85", x"0f85", x"0f85", x"0f85", x"0f85", x"0f85", x"0f85", x"0f85", x"0f85", x"0f85", x"0f86", x"0f86", x"0f86", x"0f86", x"0f86", x"0f86", x"0f86", x"0f86", x"0f86", x"0f86", x"0f86", x"0f86", x"0f86", x"0f86", x"0f86", x"0f86", x"0f86", x"0f86", x"0f86", x"0f86", x"0f86", x"0f86", x"0f86", x"0f86", x"0f86", x"0f86", x"0f86", x"0f86", x"0f86", x"0f86", x"0f86", x"0f86", x"0f86", x"0f86", x"0f86", x"0f87", x"0f87", x"0f87", x"0f87", x"0f87", x"0f87", x"0f87", x"0f87", x"0f87", x"0f87", x"0f87", x"0f87", x"0f87", x"0f87", x"0f87", x"0f87", x"0f87", x"0f87", x"0f87", x"0f87", x"0f87", x"0f87", x"0f87", x"0f87", x"0f87", x"0f87", x"0f87", x"0f87", x"0f87", x"0f87", x"0f87", x"0f87", x"0f87", x"0f87", x"0f87", x"0f88", x"0f88", x"0f88", x"0f88", x"0f88", x"0f88", x"0f88", x"0f88", x"0f88", x"0f88", x"0f88", x"0f88", x"0f88", x"0f88", x"0f88", x"0f88", x"0f88", x"0f88", x"0f88", x"0f88", x"0f88", x"0f88", x"0f88", x"0f88", x"0f88", x"0f88", x"0f88", x"0f88", x"0f88", x"0f88", x"0f88", x"0f88", x"0f88", x"0f88", x"0f88", x"0f88", x"0f89", x"0f89", x"0f89", x"0f89", x"0f89", x"0f89", x"0f89", x"0f89", x"0f89", x"0f89", x"0f89", x"0f89", x"0f89", x"0f89", x"0f89", x"0f89", x"0f89", x"0f89", x"0f89", x"0f89", x"0f89", x"0f89", x"0f89", x"0f89", x"0f89", x"0f89", x"0f89", x"0f89", x"0f89", x"0f89", x"0f89", x"0f89", x"0f89", x"0f89", x"0f89", x"0f8a", x"0f8a", x"0f8a", x"0f8a", x"0f8a", x"0f8a", x"0f8a", x"0f8a", x"0f8a", x"0f8a", x"0f8a", x"0f8a", x"0f8a", x"0f8a", x"0f8a", x"0f8a", x"0f8a", x"0f8a", x"0f8a", x"0f8a", x"0f8a", x"0f8a", x"0f8a", x"0f8a", x"0f8a", x"0f8a", x"0f8a", x"0f8a", x"0f8a", x"0f8a", x"0f8a", x"0f8a", x"0f8a", x"0f8a", x"0f8a", x"0f8a", x"0f8a", x"0f8b", x"0f8b", x"0f8b", x"0f8b", x"0f8b", x"0f8b", x"0f8b", x"0f8b", x"0f8b", x"0f8b", x"0f8b", x"0f8b", x"0f8b", x"0f8b", x"0f8b", x"0f8b", x"0f8b", x"0f8b", x"0f8b", x"0f8b", x"0f8b", x"0f8b", x"0f8b", x"0f8b", x"0f8b", x"0f8b", x"0f8b", x"0f8b", x"0f8b", x"0f8b", x"0f8b", x"0f8b", x"0f8b", x"0f8b", x"0f8b", x"0f8b", x"0f8c", x"0f8c", x"0f8c", x"0f8c", x"0f8c", x"0f8c", x"0f8c", x"0f8c", x"0f8c", x"0f8c", x"0f8c", x"0f8c", x"0f8c", x"0f8c", x"0f8c", x"0f8c", x"0f8c", x"0f8c", x"0f8c", x"0f8c", x"0f8c", x"0f8c", x"0f8c", x"0f8c", x"0f8c", x"0f8c", x"0f8c", x"0f8c", x"0f8c", x"0f8c", x"0f8c", x"0f8c", x"0f8c", x"0f8c", x"0f8c", x"0f8c", x"0f8c", x"0f8d", x"0f8d", x"0f8d", x"0f8d", x"0f8d", x"0f8d", x"0f8d", x"0f8d", x"0f8d", x"0f8d", x"0f8d", x"0f8d", x"0f8d", x"0f8d", x"0f8d", x"0f8d", x"0f8d", x"0f8d", x"0f8d", x"0f8d", x"0f8d", x"0f8d", x"0f8d", x"0f8d", x"0f8d", x"0f8d", x"0f8d", x"0f8d", x"0f8d", x"0f8d", x"0f8d", x"0f8d", x"0f8d", x"0f8d", x"0f8d", x"0f8d", x"0f8d", x"0f8e", x"0f8e", x"0f8e", x"0f8e", x"0f8e", x"0f8e", x"0f8e", x"0f8e", x"0f8e", x"0f8e", x"0f8e", x"0f8e", x"0f8e", x"0f8e", x"0f8e", x"0f8e", x"0f8e", x"0f8e", x"0f8e", x"0f8e", x"0f8e", x"0f8e", x"0f8e", x"0f8e", x"0f8e", x"0f8e", x"0f8e", x"0f8e", x"0f8e", x"0f8e", x"0f8e", x"0f8e", x"0f8e", x"0f8e", x"0f8e", x"0f8e", x"0f8e", x"0f8e", x"0f8f", x"0f8f", x"0f8f", x"0f8f", x"0f8f", x"0f8f", x"0f8f", x"0f8f", x"0f8f", x"0f8f", x"0f8f", x"0f8f", x"0f8f", x"0f8f", x"0f8f", x"0f8f", x"0f8f", x"0f8f", x"0f8f", x"0f8f", x"0f8f", x"0f8f", x"0f8f", x"0f8f", x"0f8f", x"0f8f", x"0f8f", x"0f8f", x"0f8f", x"0f8f", x"0f8f", x"0f8f", x"0f8f", x"0f8f", x"0f8f", x"0f8f", x"0f8f", x"0f90", x"0f90", x"0f90", x"0f90", x"0f90", x"0f90", x"0f90", x"0f90", x"0f90", x"0f90", x"0f90", x"0f90", x"0f90", x"0f90", x"0f90", x"0f90", x"0f90", x"0f90", x"0f90", x"0f90", x"0f90", x"0f90", x"0f90", x"0f90", x"0f90", x"0f90", x"0f90", x"0f90", x"0f90", x"0f90", x"0f90", x"0f90", x"0f90", x"0f90", x"0f90", x"0f90", x"0f90", x"0f90", x"0f91", x"0f91", x"0f91", x"0f91", x"0f91", x"0f91", x"0f91", x"0f91", x"0f91", x"0f91", x"0f91", x"0f91", x"0f91", x"0f91", x"0f91", x"0f91", x"0f91", x"0f91", x"0f91", x"0f91", x"0f91", x"0f91", x"0f91", x"0f91", x"0f91", x"0f91", x"0f91", x"0f91", x"0f91", x"0f91", x"0f91", x"0f91", x"0f91", x"0f91", x"0f91", x"0f91", x"0f91", x"0f91", x"0f91", x"0f92", x"0f92", x"0f92", x"0f92", x"0f92", x"0f92", x"0f92", x"0f92", x"0f92", x"0f92", x"0f92", x"0f92", x"0f92", x"0f92", x"0f92", x"0f92", x"0f92", x"0f92", x"0f92", x"0f92", x"0f92", x"0f92", x"0f92", x"0f92", x"0f92", x"0f92", x"0f92", x"0f92", x"0f92", x"0f92", x"0f92", x"0f92", x"0f92", x"0f92", x"0f92", x"0f92", x"0f92", x"0f92", x"0f92", x"0f93", x"0f93", x"0f93", x"0f93", x"0f93", x"0f93", x"0f93", x"0f93", x"0f93", x"0f93", x"0f93", x"0f93", x"0f93", x"0f93", x"0f93", x"0f93", x"0f93", x"0f93", x"0f93", x"0f93", x"0f93", x"0f93", x"0f93", x"0f93", x"0f93", x"0f93", x"0f93", x"0f93", x"0f93", x"0f93", x"0f93", x"0f93", x"0f93", x"0f93", x"0f93", x"0f93", x"0f93", x"0f93", x"0f93", x"0f94", x"0f94", x"0f94", x"0f94", x"0f94", x"0f94", x"0f94", x"0f94", x"0f94", x"0f94", x"0f94", x"0f94", x"0f94", x"0f94", x"0f94", x"0f94", x"0f94", x"0f94", x"0f94", x"0f94", x"0f94", x"0f94", x"0f94", x"0f94", x"0f94", x"0f94", x"0f94", x"0f94", x"0f94", x"0f94", x"0f94", x"0f94", x"0f94", x"0f94", x"0f94", x"0f94", x"0f94", x"0f94", x"0f94", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f95", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f96", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f97", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f98", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f99", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9a", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9b", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9c", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9d", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9e", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0f9f", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa0", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa1", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa2", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa3", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa4", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa5", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa6", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa7", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa8", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0fa9", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0faa", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fab", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fac", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fad", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0fae", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0faf", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb0", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb1", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb2", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb3", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb4", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb5", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb6", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb7", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb8", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fb9", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fba", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbb", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbc", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbd", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbe", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fbf", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc0", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc1", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc2", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc3", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc4", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc5", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc6", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc7", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc8", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fc9", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fca", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcb", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcc", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fcd", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fce", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fcf", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd0", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd1", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd2", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd3", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd4", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd5", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd6", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd7", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd8", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fd9", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fda", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdb", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdc", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fdd", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fde", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fdf", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe0", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe1", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe2", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe3", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe4", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe5", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe6", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe7", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe8", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fe9", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0fea", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0feb", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fec", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fed", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fee", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0fef", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff0", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff1", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff2", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff3", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff4", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff5", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff6", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff7", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff8", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ff9", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffa", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffb", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffc", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0ffd", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0002", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0003", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0004", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0005", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0006", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0007", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0008", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"0009", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000a", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000b", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000c", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000d", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000e", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"000f", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0010", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0011", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0012", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0013", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0014", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0015", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0016", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0017", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0018", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"0019", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001a", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001b", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001c", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001d", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001e", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"001f", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0020", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0021", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0022", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0023", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0024", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0025", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0026", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0027", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0028", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"0029", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002a", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002b", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002c", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002d", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002e", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"002f", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0030", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0031", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0032", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0033", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0034", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0035", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0036", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0037", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0038", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"0039", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003a", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003b", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003c", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003d", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003e", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"003f", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0040", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0041", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0042", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0043", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0044", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0045", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0046", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0047", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0048", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"0049", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004a", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004b", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004c", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004d", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004e", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"004f", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0050", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0051", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0052", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0053", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0054", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0055", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0056", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0057", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0058", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"0059", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005a", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005b", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005c", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005d", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005e", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"005f", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0060", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0061", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0062", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0063", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0064", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0065", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0066", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0067", x"0068", x"0068", x"0068", x"0068", x"0068", x"0068", x"0068", x"0068", x"0068", x"0068", x"0068", x"0068", x"0068", x"0068", x"0068", x"0068", x"0068", x"0068", x"0068", x"0068", x"0068", x"0068", x"0068", x"0068", x"0068", x"0068", x"0068", x"0068", x"0068", x"0068", x"0068", x"0068", x"0068", x"0068", x"0068", x"0068", x"0068", x"0068", x"0068", x"0068", x"0069", x"0069", x"0069", x"0069", x"0069", x"0069", x"0069", x"0069", x"0069", x"0069", x"0069", x"0069", x"0069", x"0069", x"0069", x"0069", x"0069", x"0069", x"0069", x"0069", x"0069", x"0069", x"0069", x"0069", x"0069", x"0069", x"0069", x"0069", x"0069", x"0069", x"0069", x"0069", x"0069", x"0069", x"0069", x"0069", x"0069", x"0069", x"0069", x"0069", x"006a", x"006a", x"006a", x"006a", x"006a", x"006a", x"006a", x"006a", x"006a", x"006a", x"006a", x"006a", x"006a", x"006a", x"006a", x"006a", x"006a", x"006a", x"006a", x"006a", x"006a", x"006a", x"006a", x"006a", x"006a", x"006a", x"006a", x"006a", x"006a", x"006a", x"006a", x"006a", x"006a", x"006a", x"006a", x"006a", x"006a", x"006a", x"006a", x"006b", x"006b", x"006b", x"006b", x"006b", x"006b", x"006b", x"006b", x"006b", x"006b", x"006b", x"006b", x"006b", x"006b", x"006b", x"006b", x"006b", x"006b", x"006b", x"006b", x"006b", x"006b", x"006b", x"006b", x"006b", x"006b", x"006b", x"006b", x"006b", x"006b", x"006b", x"006b", x"006b", x"006b", x"006b", x"006b", x"006b", x"006b", x"006b", x"006c", x"006c", x"006c", x"006c", x"006c", x"006c", x"006c", x"006c", x"006c", x"006c", x"006c", x"006c", x"006c", x"006c", x"006c", x"006c", x"006c", x"006c", x"006c", x"006c", x"006c", x"006c", x"006c", x"006c", x"006c", x"006c", x"006c", x"006c", x"006c", x"006c", x"006c", x"006c", x"006c", x"006c", x"006c", x"006c", x"006c", x"006c", x"006c", x"006d", x"006d", x"006d", x"006d", x"006d", x"006d", x"006d", x"006d", x"006d", x"006d", x"006d", x"006d", x"006d", x"006d", x"006d", x"006d", x"006d", x"006d", x"006d", x"006d", x"006d", x"006d", x"006d", x"006d", x"006d", x"006d", x"006d", x"006d", x"006d", x"006d", x"006d", x"006d", x"006d", x"006d", x"006d", x"006d", x"006d", x"006d", x"006d", x"006e", x"006e", x"006e", x"006e", x"006e", x"006e", x"006e", x"006e", x"006e", x"006e", x"006e", x"006e", x"006e", x"006e", x"006e", x"006e", x"006e", x"006e", x"006e", x"006e", x"006e", x"006e", x"006e", x"006e", x"006e", x"006e", x"006e", x"006e", x"006e", x"006e", x"006e", x"006e", x"006e", x"006e", x"006e", x"006e", x"006e", x"006e", x"006f", x"006f", x"006f", x"006f", x"006f", x"006f", x"006f", x"006f", x"006f", x"006f", x"006f", x"006f", x"006f", x"006f", x"006f", x"006f", x"006f", x"006f", x"006f", x"006f", x"006f", x"006f", x"006f", x"006f", x"006f", x"006f", x"006f", x"006f", x"006f", x"006f", x"006f", x"006f", x"006f", x"006f", x"006f", x"006f", x"006f", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0070", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0071", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0072", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0073", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0074", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0075", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0076", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0077", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0078", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"0079", x"007a", x"007a", x"007a", x"007a", x"007a", x"007a", x"007a", x"007a", x"007a", x"007a", x"007a", x"007a", x"007a", x"007a", x"007a", x"007a", x"007a", x"007a", x"007a", x"007a", x"007a", x"007a", x"007a", x"007a", x"007a", x"007a", x"007a", x"007a", x"007a", x"007a", x"007a", x"007a", x"007a", x"007a", x"007a", x"007b", x"007b", x"007b", x"007b", x"007b", x"007b", x"007b", x"007b", x"007b", x"007b", x"007b", x"007b", x"007b", x"007b", x"007b", x"007b", x"007b", x"007b", x"007b", x"007b", x"007b", x"007b", x"007b", x"007b", x"007b", x"007b", x"007b", x"007b", x"007b", x"007b", x"007b", x"007b", x"007b", x"007b", x"007c", x"007c", x"007c", x"007c", x"007c", x"007c", x"007c", x"007c", x"007c", x"007c", x"007c", x"007c", x"007c", x"007c", x"007c", x"007c", x"007c", x"007c", x"007c", x"007c", x"007c", x"007c", x"007c", x"007c", x"007c", x"007c", x"007c", x"007c", x"007c", x"007c", x"007c", x"007c", x"007c", x"007c", x"007d", x"007d", x"007d", x"007d", x"007d", x"007d", x"007d", x"007d", x"007d", x"007d", x"007d", x"007d", x"007d", x"007d", x"007d", x"007d", x"007d", x"007d", x"007d", x"007d", x"007d", x"007d", x"007d", x"007d", x"007d", x"007d", x"007d", x"007d", x"007d", x"007d", x"007d", x"007d", x"007d", x"007e", x"007e", x"007e", x"007e", x"007e", x"007e", x"007e", x"007e", x"007e", x"007e", x"007e", x"007e", x"007e", x"007e", x"007e", x"007e", x"007e", x"007e", x"007e", x"007e", x"007e", x"007e", x"007e", x"007e", x"007e", x"007e", x"007e", x"007e", x"007e", x"007e", x"007e", x"007e", x"007e", x"007e", x"007f", x"007f", x"007f", x"007f", x"007f", x"007f", x"007f", x"007f", x"007f", x"007f", x"007f", x"007f", x"007f", x"007f", x"007f", x"007f", x"007f", x"007f", x"007f", x"007f", x"007f", x"007f", x"007f", x"007f", x"007f", x"007f", x"007f", x"007f", x"007f", x"007f", x"007f", x"007f", x"007f", x"0080", x"0080", x"0080", x"0080", x"0080", x"0080", x"0080", x"0080", x"0080", x"0080", x"0080", x"0080", x"0080", x"0080", x"0080", x"0080", x"0080", x"0080", x"0080", x"0080", x"0080", x"0080", x"0080", x"0080", x"0080", x"0080", x"0080", x"0080", x"0080", x"0080", x"0080", x"0080", x"0080", x"0081", x"0081", x"0081", x"0081", x"0081", x"0081", x"0081", x"0081", x"0081", x"0081", x"0081", x"0081", x"0081", x"0081", x"0081", x"0081", x"0081", x"0081", x"0081", x"0081", x"0081", x"0081", x"0081", x"0081", x"0081", x"0081", x"0081", x"0081", x"0081", x"0081", x"0081", x"0081", x"0082", x"0082", x"0082", x"0082", x"0082", x"0082", x"0082", x"0082", x"0082", x"0082", x"0082", x"0082", x"0082", x"0082", x"0082", x"0082", x"0082", x"0082", x"0082", x"0082", x"0082", x"0082", x"0082", x"0082", x"0082", x"0082", x"0082", x"0082", x"0082", x"0082", x"0082", x"0082", x"0082", x"0083", x"0083", x"0083", x"0083", x"0083", x"0083", x"0083", x"0083", x"0083", x"0083", x"0083", x"0083", x"0083", x"0083", x"0083", x"0083", x"0083", x"0083", x"0083", x"0083", x"0083", x"0083", x"0083", x"0083", x"0083", x"0083", x"0083", x"0083", x"0083", x"0083", x"0083", x"0083", x"0084", x"0084", x"0084", x"0084", x"0084", x"0084", x"0084", x"0084", x"0084", x"0084", x"0084", x"0084", x"0084", x"0084", x"0084", x"0084", x"0084", x"0084", x"0084", x"0084", x"0084", x"0084", x"0084", x"0084", x"0084", x"0084", x"0084", x"0084", x"0084", x"0084", x"0084", x"0084", x"0085", x"0085", x"0085", x"0085", x"0085", x"0085", x"0085", x"0085", x"0085", x"0085", x"0085", x"0085", x"0085", x"0085", x"0085", x"0085", x"0085", x"0085", x"0085", x"0085", x"0085", x"0085", x"0085", x"0085", x"0085", x"0085", x"0085", x"0085", x"0085", x"0085", x"0085", x"0085", x"0086", x"0086", x"0086", x"0086", x"0086", x"0086", x"0086", x"0086", x"0086", x"0086", x"0086", x"0086", x"0086", x"0086", x"0086", x"0086", x"0086", x"0086", x"0086", x"0086", x"0086", x"0086", x"0086", x"0086", x"0086", x"0086", x"0086", x"0086", x"0086", x"0086", x"0086", x"0087", x"0087", x"0087", x"0087", x"0087", x"0087", x"0087", x"0087", x"0087", x"0087", x"0087", x"0087", x"0087", x"0087", x"0087", x"0087", x"0087", x"0087", x"0087", x"0087", x"0087", x"0087", x"0087", x"0087", x"0087", x"0087", x"0087", x"0087", x"0087", x"0087", x"0087", x"0087", x"0088", x"0088", x"0088", x"0088", x"0088", x"0088", x"0088", x"0088", x"0088", x"0088", x"0088", x"0088", x"0088", x"0088", x"0088", x"0088", x"0088", x"0088", x"0088", x"0088", x"0088", x"0088", x"0088", x"0088", x"0088", x"0088", x"0088", x"0088", x"0088", x"0088", x"0088", x"0089", x"0089", x"0089", x"0089", x"0089", x"0089", x"0089", x"0089", x"0089", x"0089", x"0089", x"0089", x"0089", x"0089", x"0089", x"0089", x"0089", x"0089", x"0089", x"0089", x"0089", x"0089", x"0089", x"0089", x"0089", x"0089", x"0089", x"0089", x"0089", x"0089", x"008a", x"008a", x"008a", x"008a", x"008a", x"008a", x"008a", x"008a", x"008a", x"008a", x"008a", x"008a", x"008a", x"008a", x"008a", x"008a", x"008a", x"008a", x"008a", x"008a", x"008a", x"008a", x"008a", x"008a", x"008a", x"008a", x"008a", x"008a", x"008a", x"008a", x"008a", x"008b", x"008b", x"008b", x"008b", x"008b", x"008b", x"008b", x"008b", x"008b", x"008b", x"008b", x"008b", x"008b", x"008b", x"008b", x"008b", x"008b", x"008b", x"008b", x"008b", x"008b", x"008b", x"008b", x"008b", x"008b", x"008b", x"008b", x"008b", x"008b", x"008b", x"008c", x"008c", x"008c", x"008c", x"008c", x"008c", x"008c", x"008c", x"008c", x"008c", x"008c", x"008c", x"008c", x"008c", x"008c", x"008c", x"008c", x"008c", x"008c", x"008c", x"008c", x"008c", x"008c", x"008c", x"008c", x"008c", x"008c", x"008c", x"008c", x"008c", x"008c", x"008d", x"008d", x"008d", x"008d", x"008d", x"008d", x"008d", x"008d", x"008d", x"008d", x"008d", x"008d", x"008d", x"008d", x"008d", x"008d", x"008d", x"008d", x"008d", x"008d", x"008d", x"008d", x"008d", x"008d", x"008d", x"008d", x"008d", x"008d", x"008d", x"008d", x"008e", x"008e", x"008e", x"008e", x"008e", x"008e", x"008e", x"008e", x"008e", x"008e", x"008e", x"008e", x"008e", x"008e", x"008e", x"008e", x"008e", x"008e", x"008e", x"008e", x"008e", x"008e", x"008e", x"008e", x"008e", x"008e", x"008e", x"008e", x"008e", x"008f", x"008f", x"008f", x"008f", x"008f", x"008f", x"008f", x"008f", x"008f", x"008f", x"008f", x"008f", x"008f", x"008f", x"008f", x"008f", x"008f", x"008f", x"008f", x"008f", x"008f", x"008f", x"008f", x"008f", x"008f", x"008f", x"008f", x"008f", x"008f", x"008f", x"0090", x"0090", x"0090", x"0090", x"0090", x"0090", x"0090", x"0090", x"0090", x"0090", x"0090", x"0090", x"0090", x"0090", x"0090", x"0090", x"0090", x"0090", x"0090", x"0090", x"0090", x"0090", x"0090", x"0090", x"0090", x"0090", x"0090", x"0090", x"0090", x"0091", x"0091", x"0091", x"0091", x"0091", x"0091", x"0091", x"0091", x"0091", x"0091", x"0091", x"0091", x"0091", x"0091", x"0091", x"0091", x"0091", x"0091", x"0091", x"0091", x"0091", x"0091", x"0091", x"0091", x"0091", x"0091", x"0091", x"0091", x"0091", x"0092", x"0092", x"0092", x"0092", x"0092", x"0092", x"0092", x"0092", x"0092", x"0092", x"0092", x"0092", x"0092", x"0092", x"0092", x"0092", x"0092", x"0092", x"0092", x"0092", x"0092", x"0092", x"0092", x"0092", x"0092", x"0092", x"0092", x"0092", x"0092", x"0093", x"0093", x"0093", x"0093", x"0093", x"0093", x"0093", x"0093", x"0093", x"0093", x"0093", x"0093", x"0093", x"0093", x"0093", x"0093", x"0093", x"0093", x"0093", x"0093", x"0093", x"0093", x"0093", x"0093", x"0093", x"0093", x"0093", x"0093", x"0093", x"0094", x"0094", x"0094", x"0094", x"0094", x"0094", x"0094", x"0094", x"0094", x"0094", x"0094", x"0094", x"0094", x"0094", x"0094", x"0094", x"0094", x"0094", x"0094", x"0094", x"0094", x"0094", x"0094", x"0094", x"0094", x"0094", x"0094", x"0094", x"0094", x"0095", x"0095", x"0095", x"0095", x"0095", x"0095", x"0095", x"0095", x"0095", x"0095", x"0095", x"0095", x"0095", x"0095", x"0095", x"0095", x"0095", x"0095", x"0095", x"0095", x"0095", x"0095", x"0095", x"0095", x"0095", x"0095", x"0095", x"0095", x"0096", x"0096", x"0096", x"0096", x"0096", x"0096", x"0096", x"0096", x"0096", x"0096", x"0096", x"0096", x"0096", x"0096", x"0096", x"0096", x"0096", x"0096", x"0096", x"0096", x"0096", x"0096", x"0096", x"0096", x"0096", x"0096", x"0096", x"0096", x"0096", x"0097", x"0097", x"0097", x"0097", x"0097", x"0097", x"0097", x"0097", x"0097", x"0097", x"0097", x"0097", x"0097", x"0097", x"0097", x"0097", x"0097", x"0097", x"0097", x"0097", x"0097", x"0097", x"0097", x"0097", x"0097", x"0097", x"0097", x"0097", x"0098", x"0098", x"0098", x"0098", x"0098", x"0098", x"0098", x"0098", x"0098", x"0098", x"0098", x"0098", x"0098", x"0098", x"0098", x"0098", x"0098", x"0098", x"0098", x"0098", x"0098", x"0098", x"0098", x"0098", x"0098", x"0098", x"0098", x"0098", x"0099", x"0099", x"0099", x"0099", x"0099", x"0099", x"0099", x"0099", x"0099", x"0099", x"0099", x"0099", x"0099", x"0099", x"0099", x"0099", x"0099", x"0099", x"0099", x"0099", x"0099", x"0099", x"0099", x"0099", x"0099", x"0099", x"0099", x"009a", x"009a", x"009a", x"009a", x"009a", x"009a", x"009a", x"009a", x"009a", x"009a", x"009a", x"009a", x"009a", x"009a", x"009a", x"009a", x"009a", x"009a", x"009a", x"009a", x"009a", x"009a", x"009a", x"009a", x"009a", x"009a", x"009a", x"009a", x"009b", x"009b", x"009b", x"009b", x"009b", x"009b", x"009b", x"009b", x"009b", x"009b", x"009b", x"009b", x"009b", x"009b", x"009b", x"009b", x"009b", x"009b", x"009b", x"009b", x"009b", x"009b", x"009b", x"009b", x"009b", x"009b", x"009b", x"009c", x"009c", x"009c", x"009c", x"009c", x"009c", x"009c", x"009c", x"009c", x"009c", x"009c", x"009c", x"009c", x"009c", x"009c", x"009c", x"009c", x"009c", x"009c", x"009c", x"009c", x"009c", x"009c", x"009c", x"009c", x"009c", x"009c", x"009d", x"009d", x"009d", x"009d", x"009d", x"009d", x"009d", x"009d", x"009d", x"009d", x"009d", x"009d", x"009d", x"009d", x"009d", x"009d", x"009d", x"009d", x"009d", x"009d", x"009d", x"009d", x"009d", x"009d", x"009d", x"009d", x"009d", x"009e", x"009e", x"009e", x"009e", x"009e", x"009e", x"009e", x"009e", x"009e", x"009e", x"009e", x"009e", x"009e", x"009e", x"009e", x"009e", x"009e", x"009e", x"009e", x"009e", x"009e", x"009e", x"009e", x"009e", x"009e", x"009e", x"009e", x"009f", x"009f", x"009f", x"009f", x"009f", x"009f", x"009f", x"009f", x"009f", x"009f", x"009f", x"009f", x"009f", x"009f", x"009f", x"009f", x"009f", x"009f", x"009f", x"009f", x"009f", x"009f", x"009f", x"009f", x"009f", x"009f", x"009f", x"00a0", x"00a0", x"00a0", x"00a0", x"00a0", x"00a0", x"00a0", x"00a0", x"00a0", x"00a0", x"00a0", x"00a0", x"00a0", x"00a0", x"00a0", x"00a0", x"00a0", x"00a0", x"00a0", x"00a0", x"00a0", x"00a0", x"00a0", x"00a0", x"00a0", x"00a0", x"00a0", x"00a1", x"00a1", x"00a1", x"00a1", x"00a1", x"00a1", x"00a1", x"00a1", x"00a1", x"00a1", x"00a1", x"00a1", x"00a1", x"00a1", x"00a1", x"00a1", x"00a1", x"00a1", x"00a1", x"00a1", x"00a1", x"00a1", x"00a1", x"00a1", x"00a1", x"00a1", x"00a2", x"00a2", x"00a2", x"00a2", x"00a2", x"00a2", x"00a2", x"00a2", x"00a2", x"00a2", x"00a2", x"00a2", x"00a2", x"00a2", x"00a2", x"00a2", x"00a2", x"00a2", x"00a2", x"00a2", x"00a2", x"00a2", x"00a2", x"00a2", x"00a2", x"00a2", x"00a3", x"00a3", x"00a3", x"00a3", x"00a3", x"00a3", x"00a3", x"00a3", x"00a3", x"00a3", x"00a3", x"00a3", x"00a3", x"00a3", x"00a3", x"00a3", x"00a3", x"00a3", x"00a3", x"00a3", x"00a3", x"00a3", x"00a3", x"00a3", x"00a3", x"00a3", x"00a4", x"00a4", x"00a4", x"00a4", x"00a4", x"00a4", x"00a4", x"00a4", x"00a4", x"00a4", x"00a4", x"00a4", x"00a4", x"00a4", x"00a4", x"00a4", x"00a4", x"00a4", x"00a4", x"00a4", x"00a4", x"00a4", x"00a4", x"00a4", x"00a4", x"00a4", x"00a5", x"00a5", x"00a5", x"00a5", x"00a5", x"00a5", x"00a5", x"00a5", x"00a5", x"00a5", x"00a5", x"00a5", x"00a5", x"00a5", x"00a5", x"00a5", x"00a5", x"00a5", x"00a5", x"00a5", x"00a5", x"00a5", x"00a5", x"00a5", x"00a5", x"00a5", x"00a6", x"00a6", x"00a6", x"00a6", x"00a6", x"00a6", x"00a6", x"00a6", x"00a6", x"00a6", x"00a6", x"00a6", x"00a6", x"00a6", x"00a6", x"00a6", x"00a6", x"00a6", x"00a6", x"00a6", x"00a6", x"00a6", x"00a6", x"00a6", x"00a6", x"00a6", x"00a7", x"00a7", x"00a7", x"00a7", x"00a7", x"00a7", x"00a7", x"00a7", x"00a7", x"00a7", x"00a7", x"00a7", x"00a7", x"00a7", x"00a7", x"00a7", x"00a7", x"00a7", x"00a7", x"00a7", x"00a7", x"00a7", x"00a7", x"00a7", x"00a7", x"00a8", x"00a8", x"00a8", x"00a8", x"00a8", x"00a8", x"00a8", x"00a8", x"00a8", x"00a8", x"00a8", x"00a8", x"00a8", x"00a8", x"00a8", x"00a8", x"00a8", x"00a8", x"00a8", x"00a8", x"00a8", x"00a8", x"00a8", x"00a8", x"00a8", x"00a8", x"00a9", x"00a9", x"00a9", x"00a9", x"00a9", x"00a9", x"00a9", x"00a9", x"00a9", x"00a9", x"00a9", x"00a9", x"00a9", x"00a9", x"00a9", x"00a9", x"00a9", x"00a9", x"00a9", x"00a9", x"00a9", x"00a9", x"00a9", x"00a9", x"00a9", x"00aa", x"00aa", x"00aa", x"00aa", x"00aa", x"00aa", x"00aa", x"00aa", x"00aa", x"00aa", x"00aa", x"00aa", x"00aa", x"00aa", x"00aa", x"00aa", x"00aa", x"00aa", x"00aa", x"00aa", x"00aa", x"00aa", x"00aa", x"00aa", x"00aa", x"00ab", x"00ab", x"00ab", x"00ab", x"00ab", x"00ab", x"00ab", x"00ab", x"00ab", x"00ab", x"00ab", x"00ab", x"00ab", x"00ab", x"00ab", x"00ab", x"00ab", x"00ab", x"00ab", x"00ab", x"00ab", x"00ab", x"00ab", x"00ab", x"00ab", x"00ac", x"00ac", x"00ac", x"00ac", x"00ac", x"00ac", x"00ac", x"00ac", x"00ac", x"00ac", x"00ac", x"00ac", x"00ac", x"00ac", x"00ac", x"00ac", x"00ac", x"00ac", x"00ac", x"00ac", x"00ac", x"00ac", x"00ac", x"00ac", x"00ac", x"00ad", x"00ad", x"00ad", x"00ad", x"00ad", x"00ad", x"00ad", x"00ad", x"00ad", x"00ad", x"00ad", x"00ad", x"00ad", x"00ad", x"00ad", x"00ad", x"00ad", x"00ad", x"00ad", x"00ad", x"00ad", x"00ad", x"00ad", x"00ad", x"00ae", x"00ae", x"00ae", x"00ae", x"00ae", x"00ae", x"00ae", x"00ae", x"00ae", x"00ae", x"00ae", x"00ae", x"00ae", x"00ae", x"00ae", x"00ae", x"00ae", x"00ae", x"00ae", x"00ae", x"00ae", x"00ae", x"00ae", x"00ae", x"00ae", x"00af", x"00af", x"00af", x"00af", x"00af", x"00af", x"00af", x"00af", x"00af", x"00af", x"00af", x"00af", x"00af", x"00af", x"00af", x"00af", x"00af", x"00af", x"00af", x"00af", x"00af", x"00af", x"00af", x"00af", x"00b0", x"00b0", x"00b0", x"00b0", x"00b0", x"00b0", x"00b0", x"00b0", x"00b0", x"00b0", x"00b0", x"00b0", x"00b0", x"00b0", x"00b0", x"00b0", x"00b0", x"00b0", x"00b0", x"00b0", x"00b0", x"00b0", x"00b0", x"00b0", x"00b1", x"00b1", x"00b1", x"00b1", x"00b1", x"00b1", x"00b1", x"00b1", x"00b1", x"00b1", x"00b1", x"00b1", x"00b1", x"00b1", x"00b1", x"00b1", x"00b1", x"00b1", x"00b1", x"00b1", x"00b1", x"00b1", x"00b1", x"00b1", x"00b1", x"00b2", x"00b2", x"00b2", x"00b2", x"00b2", x"00b2", x"00b2", x"00b2", x"00b2", x"00b2", x"00b2", x"00b2", x"00b2", x"00b2", x"00b2", x"00b2", x"00b2", x"00b2", x"00b2", x"00b2", x"00b2", x"00b2", x"00b2", x"00b2", x"00b3", x"00b3", x"00b3", x"00b3", x"00b3", x"00b3", x"00b3", x"00b3", x"00b3", x"00b3", x"00b3", x"00b3", x"00b3", x"00b3", x"00b3", x"00b3", x"00b3", x"00b3", x"00b3", x"00b3", x"00b3", x"00b3", x"00b3", x"00b4", x"00b4", x"00b4", x"00b4", x"00b4", x"00b4", x"00b4", x"00b4", x"00b4", x"00b4", x"00b4", x"00b4", x"00b4", x"00b4", x"00b4", x"00b4", x"00b4", x"00b4", x"00b4", x"00b4", x"00b4", x"00b4", x"00b4", x"00b4", x"00b5", x"00b5", x"00b5", x"00b5", x"00b5", x"00b5", x"00b5", x"00b5", x"00b5", x"00b5", x"00b5", x"00b5", x"00b5", x"00b5", x"00b5", x"00b5", x"00b5", x"00b5", x"00b5", x"00b5", x"00b5", x"00b5", x"00b5", x"00b5", x"00b6", x"00b6", x"00b6", x"00b6", x"00b6", x"00b6", x"00b6", x"00b6", x"00b6", x"00b6", x"00b6", x"00b6", x"00b6", x"00b6", x"00b6", x"00b6", x"00b6", x"00b6", x"00b6", x"00b6", x"00b6", x"00b6", x"00b6", x"00b7", x"00b7", x"00b7", x"00b7", x"00b7", x"00b7", x"00b7", x"00b7", x"00b7", x"00b7", x"00b7", x"00b7", x"00b7", x"00b7", x"00b7", x"00b7", x"00b7", x"00b7", x"00b7", x"00b7", x"00b7", x"00b7", x"00b7", x"00b7", x"00b8", x"00b8", x"00b8", x"00b8", x"00b8", x"00b8", x"00b8", x"00b8", x"00b8", x"00b8", x"00b8", x"00b8", x"00b8", x"00b8", x"00b8", x"00b8", x"00b8", x"00b8", x"00b8", x"00b8", x"00b8", x"00b8", x"00b8", x"00b9", x"00b9", x"00b9", x"00b9", x"00b9", x"00b9", x"00b9", x"00b9", x"00b9", x"00b9", x"00b9", x"00b9", x"00b9", x"00b9", x"00b9", x"00b9", x"00b9", x"00b9", x"00b9", x"00b9", x"00b9", x"00b9", x"00b9", x"00ba", x"00ba", x"00ba", x"00ba", x"00ba", x"00ba", x"00ba", x"00ba", x"00ba", x"00ba", x"00ba", x"00ba", x"00ba", x"00ba", x"00ba", x"00ba", x"00ba", x"00ba", x"00ba", x"00ba", x"00ba", x"00ba", x"00ba", x"00bb", x"00bb", x"00bb", x"00bb", x"00bb", x"00bb", x"00bb", x"00bb", x"00bb", x"00bb", x"00bb", x"00bb", x"00bb", x"00bb", x"00bb", x"00bb", x"00bb", x"00bb", x"00bb", x"00bb", x"00bb", x"00bb", x"00bb", x"00bc", x"00bc", x"00bc", x"00bc", x"00bc", x"00bc", x"00bc", x"00bc", x"00bc", x"00bc", x"00bc", x"00bc", x"00bc", x"00bc", x"00bc", x"00bc", x"00bc", x"00bc", x"00bc", x"00bc", x"00bc", x"00bc", x"00bc", x"00bd", x"00bd", x"00bd", x"00bd", x"00bd", x"00bd", x"00bd", x"00bd", x"00bd", x"00bd", x"00bd", x"00bd", x"00bd", x"00bd", x"00bd", x"00bd", x"00bd", x"00bd", x"00bd", x"00bd", x"00bd", x"00bd", x"00be", x"00be", x"00be", x"00be", x"00be", x"00be", x"00be", x"00be", x"00be", x"00be", x"00be", x"00be", x"00be", x"00be", x"00be", x"00be", x"00be", x"00be", x"00be", x"00be", x"00be", x"00be", x"00be", x"00bf", x"00bf", x"00bf", x"00bf", x"00bf", x"00bf", x"00bf", x"00bf", x"00bf", x"00bf", x"00bf", x"00bf", x"00bf", x"00bf", x"00bf", x"00bf", x"00bf", x"00bf", x"00bf", x"00bf", x"00bf", x"00bf", x"00c0", x"00c0", x"00c0", x"00c0", x"00c0", x"00c0", x"00c0", x"00c0", x"00c0", x"00c0", x"00c0", x"00c0", x"00c0", x"00c0", x"00c0", x"00c0", x"00c0", x"00c0", x"00c0", x"00c0", x"00c0", x"00c0", x"00c0", x"00c1", x"00c1", x"00c1", x"00c1", x"00c1", x"00c1", x"00c1", x"00c1", x"00c1", x"00c1", x"00c1", x"00c1", x"00c1", x"00c1", x"00c1", x"00c1", x"00c1", x"00c1", x"00c1", x"00c1", x"00c1", x"00c1", x"00c2", x"00c2", x"00c2", x"00c2", x"00c2", x"00c2", x"00c2", x"00c2", x"00c2", x"00c2", x"00c2", x"00c2", x"00c2", x"00c2", x"00c2", x"00c2", x"00c2", x"00c2", x"00c2", x"00c2", x"00c2", x"00c2", x"00c3", x"00c3", x"00c3", x"00c3", x"00c3", x"00c3", x"00c3", x"00c3", x"00c3", x"00c3", x"00c3", x"00c3", x"00c3", x"00c3", x"00c3", x"00c3", x"00c3", x"00c3", x"00c3", x"00c3", x"00c3", x"00c3", x"00c4", x"00c4", x"00c4", x"00c4", x"00c4", x"00c4", x"00c4", x"00c4", x"00c4", x"00c4", x"00c4", x"00c4", x"00c4", x"00c4", x"00c4", x"00c4", x"00c4", x"00c4", x"00c4", x"00c4", x"00c4", x"00c4", x"00c5", x"00c5", x"00c5", x"00c5", x"00c5", x"00c5", x"00c5", x"00c5", x"00c5", x"00c5", x"00c5", x"00c5", x"00c5", x"00c5", x"00c5", x"00c5", x"00c5", x"00c5", x"00c5", x"00c5", x"00c5", x"00c5", x"00c6", x"00c6", x"00c6", x"00c6", x"00c6", x"00c6", x"00c6", x"00c6", x"00c6", x"00c6", x"00c6", x"00c6", x"00c6", x"00c6", x"00c6", x"00c6", x"00c6", x"00c6", x"00c6", x"00c6", x"00c6", x"00c7", x"00c7", x"00c7", x"00c7", x"00c7", x"00c7", x"00c7", x"00c7", x"00c7", x"00c7", x"00c7", x"00c7", x"00c7", x"00c7", x"00c7", x"00c7", x"00c7", x"00c7", x"00c7", x"00c7", x"00c7", x"00c7", x"00c8", x"00c8", x"00c8", x"00c8", x"00c8", x"00c8", x"00c8", x"00c8", x"00c8", x"00c8", x"00c8", x"00c8", x"00c8", x"00c8", x"00c8", x"00c8", x"00c8", x"00c8", x"00c8", x"00c8", x"00c8", x"00c9", x"00c9", x"00c9", x"00c9", x"00c9", x"00c9", x"00c9", x"00c9", x"00c9", x"00c9", x"00c9", x"00c9", x"00c9", x"00c9", x"00c9", x"00c9", x"00c9", x"00c9", x"00c9", x"00c9", x"00c9", x"00c9", x"00ca", x"00ca", x"00ca", x"00ca", x"00ca", x"00ca", x"00ca", x"00ca", x"00ca", x"00ca", x"00ca", x"00ca", x"00ca", x"00ca", x"00ca", x"00ca", x"00ca", x"00ca", x"00ca", x"00ca", x"00ca", x"00cb", x"00cb", x"00cb", x"00cb", x"00cb", x"00cb", x"00cb", x"00cb", x"00cb", x"00cb", x"00cb", x"00cb", x"00cb", x"00cb", x"00cb", x"00cb", x"00cb", x"00cb", x"00cb", x"00cb", x"00cb", x"00cc", x"00cc", x"00cc", x"00cc", x"00cc", x"00cc", x"00cc", x"00cc", x"00cc", x"00cc", x"00cc", x"00cc", x"00cc", x"00cc", x"00cc", x"00cc", x"00cc", x"00cc", x"00cc", x"00cc", x"00cc", x"00cd", x"00cd", x"00cd", x"00cd", x"00cd", x"00cd", x"00cd", x"00cd", x"00cd", x"00cd", x"00cd", x"00cd", x"00cd", x"00cd", x"00cd", x"00cd", x"00cd", x"00cd", x"00cd", x"00cd", x"00cd", x"00ce", x"00ce", x"00ce", x"00ce", x"00ce", x"00ce", x"00ce", x"00ce", x"00ce", x"00ce", x"00ce", x"00ce", x"00ce", x"00ce", x"00ce", x"00ce", x"00ce", x"00ce", x"00ce", x"00ce", x"00ce", x"00cf", x"00cf", x"00cf", x"00cf", x"00cf", x"00cf", x"00cf", x"00cf", x"00cf", x"00cf", x"00cf", x"00cf", x"00cf", x"00cf", x"00cf", x"00cf", x"00cf", x"00cf", x"00cf", x"00cf", x"00cf", x"00d0", x"00d0", x"00d0", x"00d0", x"00d0", x"00d0", x"00d0", x"00d0", x"00d0", x"00d0", x"00d0", x"00d0", x"00d0", x"00d0", x"00d0", x"00d0", x"00d0", x"00d0", x"00d0", x"00d0", x"00d0", x"00d1", x"00d1", x"00d1", x"00d1", x"00d1", x"00d1", x"00d1", x"00d1", x"00d1", x"00d1", x"00d1", x"00d1", x"00d1", x"00d1", x"00d1", x"00d1", x"00d1", x"00d1", x"00d1", x"00d1", x"00d2", x"00d2", x"00d2", x"00d2", x"00d2", x"00d2", x"00d2", x"00d2", x"00d2", x"00d2", x"00d2", x"00d2", x"00d2", x"00d2", x"00d2", x"00d2", x"00d2", x"00d2", x"00d2", x"00d2", x"00d2", x"00d3", x"00d3", x"00d3", x"00d3", x"00d3", x"00d3", x"00d3", x"00d3", x"00d3", x"00d3", x"00d3", x"00d3", x"00d3", x"00d3", x"00d3", x"00d3", x"00d3", x"00d3", x"00d3", x"00d3", x"00d4", x"00d4", x"00d4", x"00d4", x"00d4", x"00d4", x"00d4", x"00d4", x"00d4", x"00d4", x"00d4", x"00d4", x"00d4", x"00d4", x"00d4", x"00d4", x"00d4", x"00d4", x"00d4", x"00d4", x"00d4", x"00d5", x"00d5", x"00d5", x"00d5", x"00d5", x"00d5", x"00d5", x"00d5", x"00d5", x"00d5", x"00d5", x"00d5", x"00d5", x"00d5", x"00d5", x"00d5", x"00d5", x"00d5", x"00d5", x"00d5", x"00d6", x"00d6", x"00d6", x"00d6", x"00d6", x"00d6", x"00d6", x"00d6", x"00d6", x"00d6", x"00d6", x"00d6", x"00d6", x"00d6", x"00d6", x"00d6", x"00d6", x"00d6", x"00d6", x"00d6", x"00d7", x"00d7", x"00d7", x"00d7", x"00d7", x"00d7", x"00d7", x"00d7", x"00d7", x"00d7", x"00d7", x"00d7", x"00d7", x"00d7", x"00d7", x"00d7", x"00d7", x"00d7", x"00d7", x"00d7", x"00d8", x"00d8", x"00d8", x"00d8", x"00d8", x"00d8", x"00d8", x"00d8", x"00d8", x"00d8", x"00d8", x"00d8", x"00d8", x"00d8", x"00d8", x"00d8", x"00d8", x"00d8", x"00d8", x"00d8", x"00d9", x"00d9", x"00d9", x"00d9", x"00d9", x"00d9", x"00d9", x"00d9", x"00d9", x"00d9", x"00d9", x"00d9", x"00d9", x"00d9", x"00d9", x"00d9", x"00d9", x"00d9", x"00d9", x"00d9", x"00da", x"00da", x"00da", x"00da", x"00da", x"00da", x"00da", x"00da", x"00da", x"00da", x"00da", x"00da", x"00da", x"00da", x"00da", x"00da", x"00da", x"00da", x"00da", x"00da", x"00db", x"00db", x"00db", x"00db", x"00db", x"00db", x"00db", x"00db", x"00db", x"00db", x"00db", x"00db", x"00db", x"00db", x"00db", x"00db", x"00db", x"00db", x"00db", x"00dc", x"00dc", x"00dc", x"00dc", x"00dc", x"00dc", x"00dc", x"00dc", x"00dc", x"00dc", x"00dc", x"00dc", x"00dc", x"00dc", x"00dc", x"00dc", x"00dc", x"00dc", x"00dc", x"00dc", x"00dd", x"00dd", x"00dd", x"00dd", x"00dd", x"00dd", x"00dd", x"00dd", x"00dd", x"00dd", x"00dd", x"00dd", x"00dd", x"00dd", x"00dd", x"00dd", x"00dd", x"00dd", x"00dd", x"00dd", x"00de", x"00de", x"00de", x"00de", x"00de", x"00de", x"00de", x"00de", x"00de", x"00de", x"00de", x"00de", x"00de", x"00de", x"00de", x"00de", x"00de", x"00de", x"00de", x"00df", x"00df", x"00df", x"00df", x"00df", x"00df", x"00df", x"00df", x"00df", x"00df", x"00df", x"00df", x"00df", x"00df", x"00df", x"00df", x"00df", x"00df", x"00df", x"00e0", x"00e0", x"00e0", x"00e0", x"00e0", x"00e0", x"00e0", x"00e0", x"00e0", x"00e0", x"00e0", x"00e0", x"00e0", x"00e0", x"00e0", x"00e0", x"00e0", x"00e0", x"00e0", x"00e0", x"00e1", x"00e1", x"00e1", x"00e1", x"00e1", x"00e1", x"00e1", x"00e1", x"00e1", x"00e1", x"00e1", x"00e1", x"00e1", x"00e1", x"00e1", x"00e1", x"00e1", x"00e1", x"00e1", x"00e2", x"00e2", x"00e2", x"00e2", x"00e2", x"00e2", x"00e2", x"00e2", x"00e2", x"00e2", x"00e2", x"00e2", x"00e2", x"00e2", x"00e2", x"00e2", x"00e2", x"00e2", x"00e2", x"00e3", x"00e3", x"00e3", x"00e3", x"00e3", x"00e3", x"00e3", x"00e3", x"00e3", x"00e3", x"00e3", x"00e3", x"00e3", x"00e3", x"00e3", x"00e3", x"00e3", x"00e3", x"00e3", x"00e4", x"00e4", x"00e4", x"00e4", x"00e4", x"00e4", x"00e4", x"00e4", x"00e4", x"00e4", x"00e4", x"00e4", x"00e4", x"00e4", x"00e4", x"00e4", x"00e4", x"00e4", x"00e4", x"00e5", x"00e5", x"00e5", x"00e5", x"00e5", x"00e5", x"00e5", x"00e5", x"00e5", x"00e5", x"00e5", x"00e5", x"00e5", x"00e5", x"00e5", x"00e5", x"00e5", x"00e5", x"00e5", x"00e6", x"00e6", x"00e6", x"00e6", x"00e6", x"00e6", x"00e6", x"00e6", x"00e6", x"00e6", x"00e6", x"00e6", x"00e6", x"00e6", x"00e6", x"00e6", x"00e6", x"00e6", x"00e6", x"00e7", x"00e7", x"00e7", x"00e7", x"00e7", x"00e7", x"00e7", x"00e7", x"00e7", x"00e7", x"00e7", x"00e7", x"00e7", x"00e7", x"00e7", x"00e7", x"00e7", x"00e7", x"00e7", x"00e8", x"00e8", x"00e8", x"00e8", x"00e8", x"00e8", x"00e8", x"00e8", x"00e8", x"00e8", x"00e8", x"00e8", x"00e8", x"00e8", x"00e8", x"00e8", x"00e8", x"00e8", x"00e9", x"00e9", x"00e9", x"00e9", x"00e9", x"00e9", x"00e9", x"00e9", x"00e9", x"00e9", x"00e9", x"00e9", x"00e9", x"00e9", x"00e9", x"00e9", x"00e9", x"00e9", x"00e9", x"00ea", x"00ea", x"00ea", x"00ea", x"00ea", x"00ea", x"00ea", x"00ea", x"00ea", x"00ea", x"00ea", x"00ea", x"00ea", x"00ea", x"00ea", x"00ea", x"00ea", x"00ea", x"00eb", x"00eb", x"00eb", x"00eb", x"00eb", x"00eb", x"00eb", x"00eb", x"00eb", x"00eb", x"00eb", x"00eb", x"00eb", x"00eb", x"00eb", x"00eb", x"00eb", x"00eb", x"00eb", x"00ec", x"00ec", x"00ec", x"00ec", x"00ec", x"00ec", x"00ec", x"00ec", x"00ec", x"00ec", x"00ec", x"00ec", x"00ec", x"00ec", x"00ec", x"00ec", x"00ec", x"00ec", x"00ed", x"00ed", x"00ed", x"00ed", x"00ed", x"00ed", x"00ed", x"00ed", x"00ed", x"00ed", x"00ed", x"00ed", x"00ed", x"00ed", x"00ed", x"00ed", x"00ed", x"00ed", x"00ed", x"00ee", x"00ee", x"00ee", x"00ee", x"00ee", x"00ee", x"00ee", x"00ee", x"00ee", x"00ee", x"00ee", x"00ee", x"00ee", x"00ee", x"00ee", x"00ee", x"00ee", x"00ee", x"00ef", x"00ef", x"00ef", x"00ef", x"00ef", x"00ef", x"00ef", x"00ef", x"00ef", x"00ef", x"00ef", x"00ef", x"00ef", x"00ef", x"00ef", x"00ef", x"00ef", x"00ef", x"00f0", x"00f0", x"00f0", x"00f0", x"00f0", x"00f0", x"00f0", x"00f0", x"00f0", x"00f0", x"00f0", x"00f0", x"00f0", x"00f0", x"00f0", x"00f0", x"00f0", x"00f0", x"00f1", x"00f1", x"00f1", x"00f1", x"00f1", x"00f1", x"00f1", x"00f1", x"00f1", x"00f1", x"00f1", x"00f1", x"00f1", x"00f1", x"00f1", x"00f1", x"00f1", x"00f1", x"00f2", x"00f2", x"00f2", x"00f2", x"00f2", x"00f2", x"00f2", x"00f2", x"00f2", x"00f2", x"00f2", x"00f2", x"00f2", x"00f2", x"00f2", x"00f2", x"00f2", x"00f2", x"00f3", x"00f3", x"00f3", x"00f3", x"00f3", x"00f3", x"00f3", x"00f3", x"00f3", x"00f3", x"00f3", x"00f3", x"00f3", x"00f3", x"00f3", x"00f3", x"00f3", x"00f3", x"00f4", x"00f4", x"00f4", x"00f4", x"00f4", x"00f4", x"00f4", x"00f4", x"00f4", x"00f4", x"00f4", x"00f4", x"00f4", x"00f4", x"00f4", x"00f4", x"00f4", x"00f4", x"00f5", x"00f5", x"00f5", x"00f5", x"00f5", x"00f5", x"00f5", x"00f5", x"00f5", x"00f5", x"00f5", x"00f5", x"00f5", x"00f5", x"00f5", x"00f5", x"00f5", x"00f5", x"00f6", x"00f6", x"00f6", x"00f6", x"00f6", x"00f6", x"00f6", x"00f6", x"00f6", x"00f6", x"00f6", x"00f6", x"00f6", x"00f6", x"00f6", x"00f6", x"00f6", x"00f7", x"00f7", x"00f7", x"00f7", x"00f7", x"00f7", x"00f7", x"00f7", x"00f7", x"00f7", x"00f7", x"00f7", x"00f7", x"00f7", x"00f7", x"00f7", x"00f7", x"00f7", x"00f8", x"00f8", x"00f8", x"00f8", x"00f8", x"00f8", x"00f8", x"00f8", x"00f8", x"00f8", x"00f8", x"00f8", x"00f8", x"00f8", x"00f8", x"00f8", x"00f8", x"00f9", x"00f9", x"00f9", x"00f9", x"00f9", x"00f9", x"00f9", x"00f9", x"00f9", x"00f9", x"00f9", x"00f9", x"00f9", x"00f9", x"00f9", x"00f9", x"00f9", x"00f9", x"00fa", x"00fa", x"00fa", x"00fa", x"00fa", x"00fa", x"00fa", x"00fa", x"00fa", x"00fa", x"00fa", x"00fa", x"00fa", x"00fa", x"00fa", x"00fa", x"00fa", x"00fb", x"00fb", x"00fb", x"00fb", x"00fb", x"00fb", x"00fb", x"00fb", x"00fb", x"00fb", x"00fb", x"00fb", x"00fb", x"00fb", x"00fb", x"00fb", x"00fb", x"00fb", x"00fc", x"00fc", x"00fc", x"00fc", x"00fc", x"00fc", x"00fc", x"00fc", x"00fc", x"00fc", x"00fc", x"00fc", x"00fc", x"00fc", x"00fc", x"00fc", x"00fc", x"00fd", x"00fd", x"00fd", x"00fd", x"00fd", x"00fd", x"00fd", x"00fd", x"00fd", x"00fd", x"00fd", x"00fd", x"00fd", x"00fd", x"00fd", x"00fd", x"00fd", x"00fe", x"00fe", x"00fe", x"00fe", x"00fe", x"00fe", x"00fe", x"00fe", x"00fe", x"00fe", x"00fe", x"00fe", x"00fe", x"00fe", x"00fe", x"00fe", x"00fe", x"00ff", x"00ff", x"00ff", x"00ff", x"00ff", x"00ff", x"00ff", x"00ff", x"00ff", x"00ff", x"00ff", x"00ff", x"00ff", x"00ff", x"00ff", x"00ff", x"00ff", x"0100", x"0100", x"0100", x"0100", x"0100", x"0100", x"0100", x"0100", x"0100", x"0100", x"0100", x"0100", x"0100", x"0100", x"0100", x"0100", x"0100", x"0101", x"0101", x"0101", x"0101", x"0101", x"0101", x"0101", x"0101", x"0101", x"0101", x"0101", x"0101", x"0101", x"0101", x"0101", x"0101", x"0101", x"0102", x"0102", x"0102", x"0102", x"0102", x"0102", x"0102", x"0102", x"0102", x"0102", x"0102", x"0102", x"0102", x"0102", x"0102", x"0102", x"0102", x"0103", x"0103", x"0103", x"0103", x"0103", x"0103", x"0103", x"0103", x"0103", x"0103", x"0103", x"0103", x"0103", x"0103", x"0103", x"0103", x"0103", x"0104", x"0104", x"0104", x"0104", x"0104", x"0104", x"0104", x"0104", x"0104", x"0104", x"0104", x"0104", x"0104", x"0104", x"0104", x"0104", x"0104", x"0105", x"0105", x"0105", x"0105", x"0105", x"0105", x"0105", x"0105", x"0105", x"0105", x"0105", x"0105", x"0105", x"0105", x"0105", x"0105", x"0105", x"0106", x"0106", x"0106", x"0106", x"0106", x"0106", x"0106", x"0106", x"0106", x"0106", x"0106", x"0106", x"0106", x"0106", x"0106", x"0106", x"0107", x"0107", x"0107", x"0107", x"0107", x"0107", x"0107", x"0107", x"0107", x"0107", x"0107", x"0107", x"0107", x"0107", x"0107", x"0107", x"0107", x"0108", x"0108", x"0108", x"0108", x"0108", x"0108", x"0108", x"0108", x"0108", x"0108", x"0108", x"0108", x"0108", x"0108", x"0108", x"0108", x"0108", x"0109", x"0109", x"0109", x"0109", x"0109", x"0109", x"0109", x"0109", x"0109", x"0109", x"0109", x"0109", x"0109", x"0109", x"0109", x"0109", x"010a", x"010a", x"010a", x"010a", x"010a", x"010a", x"010a", x"010a", x"010a", x"010a", x"010a", x"010a", x"010a", x"010a", x"010a", x"010a", x"010b", x"010b", x"010b", x"010b", x"010b", x"010b", x"010b", x"010b", x"010b", x"010b", x"010b", x"010b", x"010b", x"010b", x"010b", x"010b", x"010b", x"010c", x"010c", x"010c", x"010c", x"010c", x"010c", x"010c", x"010c", x"010c", x"010c", x"010c", x"010c", x"010c", x"010c", x"010c", x"010c", x"010d", x"010d", x"010d", x"010d", x"010d", x"010d", x"010d", x"010d", x"010d", x"010d", x"010d", x"010d", x"010d", x"010d", x"010d", x"010d", x"010e", x"010e", x"010e", x"010e", x"010e", x"010e", x"010e", x"010e", x"010e", x"010e", x"010e", x"010e", x"010e", x"010e", x"010e", x"010e", x"010e", x"010f", x"010f", x"010f", x"010f", x"010f", x"010f", x"010f", x"010f", x"010f", x"010f", x"010f", x"010f", x"010f", x"010f", x"010f", x"010f", x"0110", x"0110", x"0110", x"0110", x"0110", x"0110", x"0110", x"0110", x"0110", x"0110", x"0110", x"0110", x"0110", x"0110", x"0110", x"0110", x"0111", x"0111", x"0111", x"0111", x"0111", x"0111", x"0111", x"0111", x"0111", x"0111", x"0111", x"0111", x"0111", x"0111", x"0111", x"0111", x"0112", x"0112", x"0112", x"0112", x"0112", x"0112", x"0112", x"0112", x"0112", x"0112", x"0112", x"0112", x"0112", x"0112", x"0112", x"0112", x"0113", x"0113", x"0113", x"0113", x"0113", x"0113", x"0113", x"0113", x"0113", x"0113", x"0113", x"0113", x"0113", x"0113", x"0113", x"0113", x"0114", x"0114", x"0114", x"0114", x"0114", x"0114", x"0114", x"0114", x"0114", x"0114", x"0114", x"0114", x"0114", x"0114", x"0114", x"0114", x"0115", x"0115", x"0115", x"0115", x"0115", x"0115", x"0115", x"0115", x"0115", x"0115", x"0115", x"0115", x"0115", x"0115", x"0115", x"0115", x"0116", x"0116", x"0116", x"0116", x"0116", x"0116", x"0116", x"0116", x"0116", x"0116", x"0116", x"0116", x"0116", x"0116", x"0116", x"0117", x"0117", x"0117", x"0117", x"0117", x"0117", x"0117", x"0117", x"0117", x"0117", x"0117", x"0117", x"0117", x"0117", x"0117", x"0117", x"0118", x"0118", x"0118", x"0118", x"0118", x"0118", x"0118", x"0118", x"0118", x"0118", x"0118", x"0118", x"0118", x"0118", x"0118", x"0118", x"0119", x"0119", x"0119", x"0119", x"0119", x"0119", x"0119", x"0119", x"0119", x"0119", x"0119", x"0119", x"0119", x"0119", x"0119", x"011a", x"011a", x"011a", x"011a", x"011a", x"011a", x"011a", x"011a", x"011a", x"011a", x"011a", x"011a", x"011a", x"011a", x"011a", x"011a", x"011b", x"011b", x"011b", x"011b", x"011b", x"011b", x"011b", x"011b", x"011b", x"011b", x"011b", x"011b", x"011b", x"011b", x"011b", x"011b", x"011c", x"011c", x"011c", x"011c", x"011c", x"011c", x"011c", x"011c", x"011c", x"011c", x"011c", x"011c", x"011c", x"011c", x"011c", x"011d", x"011d", x"011d", x"011d", x"011d", x"011d", x"011d", x"011d", x"011d", x"011d", x"011d", x"011d", x"011d", x"011d", x"011d", x"011e", x"011e", x"011e", x"011e", x"011e", x"011e", x"011e", x"011e", x"011e", x"011e", x"011e", x"011e", x"011e", x"011e", x"011e", x"011e", x"011f", x"011f", x"011f", x"011f", x"011f", x"011f", x"011f", x"011f", x"011f", x"011f", x"011f", x"011f", x"011f", x"011f", x"011f", x"0120", x"0120", x"0120", x"0120", x"0120", x"0120", x"0120", x"0120", x"0120", x"0120", x"0120", x"0120", x"0120", x"0120", x"0120", x"0121", x"0121", x"0121", x"0121", x"0121", x"0121", x"0121", x"0121", x"0121", x"0121", x"0121", x"0121", x"0121", x"0121", x"0121", x"0121", x"0122", x"0122", x"0122", x"0122", x"0122", x"0122", x"0122", x"0122", x"0122", x"0122", x"0122", x"0122", x"0122", x"0122", x"0122", x"0123", x"0123", x"0123", x"0123", x"0123", x"0123", x"0123", x"0123", x"0123", x"0123", x"0123", x"0123", x"0123", x"0123", x"0123", x"0124", x"0124", x"0124", x"0124", x"0124", x"0124", x"0124", x"0124", x"0124", x"0124", x"0124", x"0124", x"0124", x"0124", x"0124", x"0125", x"0125", x"0125", x"0125", x"0125", x"0125", x"0125", x"0125", x"0125", x"0125", x"0125", x"0125", x"0125", x"0125", x"0125", x"0126", x"0126", x"0126", x"0126", x"0126", x"0126", x"0126", x"0126", x"0126", x"0126", x"0126", x"0126", x"0126", x"0126", x"0126", x"0127", x"0127", x"0127", x"0127", x"0127", x"0127", x"0127", x"0127", x"0127", x"0127", x"0127", x"0127", x"0127", x"0127", x"0127", x"0128", x"0128", x"0128", x"0128", x"0128", x"0128", x"0128", x"0128", x"0128", x"0128", x"0128", x"0128", x"0128", x"0128", x"0128", x"0129", x"0129", x"0129", x"0129", x"0129", x"0129", x"0129", x"0129", x"0129", x"0129", x"0129", x"0129", x"0129", x"0129", x"0129", x"012a", x"012a", x"012a", x"012a", x"012a", x"012a", x"012a", x"012a", x"012a", x"012a", x"012a", x"012a", x"012a", x"012a", x"012a", x"012b", x"012b", x"012b", x"012b", x"012b", x"012b", x"012b", x"012b", x"012b", x"012b", x"012b", x"012b", x"012b", x"012b", x"012c", x"012c", x"012c", x"012c", x"012c", x"012c", x"012c", x"012c", x"012c", x"012c", x"012c", x"012c", x"012c", x"012c", x"012c", x"012d", x"012d", x"012d", x"012d", x"012d", x"012d", x"012d", x"012d", x"012d", x"012d", x"012d", x"012d", x"012d", x"012d", x"012d", x"012e", x"012e", x"012e", x"012e", x"012e", x"012e", x"012e", x"012e", x"012e", x"012e", x"012e", x"012e", x"012e", x"012e", x"012f", x"012f", x"012f", x"012f", x"012f", x"012f", x"012f", x"012f", x"012f", x"012f", x"012f", x"012f", x"012f", x"012f", x"012f", x"0130", x"0130", x"0130", x"0130", x"0130", x"0130", x"0130", x"0130", x"0130", x"0130", x"0130", x"0130", x"0130", x"0130", x"0131", x"0131", x"0131", x"0131", x"0131", x"0131", x"0131", x"0131", x"0131", x"0131", x"0131", x"0131", x"0131", x"0131", x"0131", x"0132", x"0132", x"0132", x"0132", x"0132", x"0132", x"0132", x"0132", x"0132", x"0132", x"0132", x"0132", x"0132", x"0132", x"0133", x"0133", x"0133", x"0133", x"0133", x"0133", x"0133", x"0133", x"0133", x"0133", x"0133", x"0133", x"0133", x"0133", x"0133", x"0134", x"0134", x"0134", x"0134", x"0134", x"0134", x"0134", x"0134", x"0134", x"0134", x"0134", x"0134", x"0134", x"0134", x"0135", x"0135", x"0135", x"0135", x"0135", x"0135", x"0135", x"0135", x"0135", x"0135", x"0135", x"0135", x"0135", x"0135", x"0136", x"0136", x"0136", x"0136", x"0136", x"0136", x"0136", x"0136", x"0136", x"0136", x"0136", x"0136", x"0136", x"0136", x"0136", x"0137", x"0137", x"0137", x"0137", x"0137", x"0137", x"0137", x"0137", x"0137", x"0137", x"0137", x"0137", x"0137", x"0137", x"0138", x"0138", x"0138", x"0138", x"0138", x"0138", x"0138", x"0138", x"0138", x"0138", x"0138", x"0138", x"0138", x"0138", x"0139", x"0139", x"0139", x"0139", x"0139", x"0139", x"0139", x"0139", x"0139", x"0139", x"0139", x"0139", x"0139", x"0139", x"013a", x"013a", x"013a", x"013a", x"013a", x"013a", x"013a", x"013a", x"013a", x"013a", x"013a", x"013a", x"013a", x"013a", x"013b", x"013b", x"013b", x"013b", x"013b", x"013b", x"013b", x"013b", x"013b", x"013b", x"013b", x"013b", x"013b", x"013b", x"013c", x"013c", x"013c", x"013c", x"013c", x"013c", x"013c", x"013c", x"013c", x"013c", x"013c", x"013c", x"013c", x"013c", x"013d", x"013d", x"013d", x"013d", x"013d", x"013d", x"013d", x"013d", x"013d", x"013d", x"013d", x"013d", x"013d", x"013d", x"013e", x"013e", x"013e", x"013e", x"013e", x"013e", x"013e", x"013e", x"013e", x"013e", x"013e", x"013e", x"013e", x"013e", x"013f", x"013f", x"013f", x"013f", x"013f", x"013f", x"013f", x"013f", x"013f", x"013f", x"013f", x"013f", x"013f", x"013f", x"0140", x"0140", x"0140", x"0140", x"0140", x"0140", x"0140", x"0140", x"0140", x"0140", x"0140", x"0140", x"0140", x"0140", x"0141", x"0141", x"0141", x"0141", x"0141", x"0141", x"0141", x"0141", x"0141", x"0141", x"0141", x"0141", x"0141", x"0141", x"0142", x"0142", x"0142", x"0142", x"0142", x"0142", x"0142", x"0142", x"0142", x"0142", x"0142", x"0142", x"0142", x"0142", x"0143", x"0143", x"0143", x"0143", x"0143", x"0143", x"0143", x"0143", x"0143", x"0143", x"0143", x"0143", x"0143", x"0144", x"0144", x"0144", x"0144", x"0144", x"0144", x"0144", x"0144", x"0144", x"0144", x"0144", x"0144", x"0144", x"0144", x"0145", x"0145", x"0145", x"0145", x"0145", x"0145", x"0145", x"0145", x"0145", x"0145", x"0145", x"0145", x"0145", x"0145", x"0146", x"0146", x"0146", x"0146", x"0146", x"0146", x"0146", x"0146", x"0146", x"0146", x"0146", x"0146", x"0146", x"0147", x"0147", x"0147", x"0147", x"0147", x"0147", x"0147", x"0147", x"0147", x"0147", x"0147", x"0147", x"0147", x"0147", x"0148", x"0148", x"0148", x"0148", x"0148", x"0148", x"0148", x"0148", x"0148", x"0148", x"0148", x"0148", x"0148", x"0148", x"0149", x"0149", x"0149", x"0149", x"0149", x"0149", x"0149", x"0149", x"0149", x"0149", x"0149", x"0149", x"0149", x"014a", x"014a", x"014a", x"014a", x"014a", x"014a", x"014a", x"014a", x"014a", x"014a", x"014a", x"014a", x"014a", x"014a", x"014b", x"014b", x"014b", x"014b", x"014b", x"014b", x"014b", x"014b", x"014b", x"014b", x"014b", x"014b", x"014b", x"014c", x"014c", x"014c", x"014c", x"014c", x"014c", x"014c", x"014c", x"014c", x"014c", x"014c", x"014c", x"014c", x"014d", x"014d", x"014d", x"014d", x"014d", x"014d", x"014d", x"014d", x"014d", x"014d", x"014d", x"014d", x"014d", x"014d", x"014e", x"014e", x"014e", x"014e", x"014e", x"014e", x"014e", x"014e", x"014e", x"014e", x"014e", x"014e", x"014e", x"014f", x"014f", x"014f", x"014f", x"014f", x"014f", x"014f", x"014f", x"014f", x"014f", x"014f", x"014f", x"014f", x"0150", x"0150", x"0150", x"0150", x"0150", x"0150", x"0150", x"0150", x"0150", x"0150", x"0150", x"0150", x"0150", x"0150", x"0151", x"0151", x"0151", x"0151", x"0151", x"0151", x"0151", x"0151", x"0151", x"0151", x"0151", x"0151", x"0151", x"0152", x"0152", x"0152", x"0152", x"0152", x"0152", x"0152", x"0152", x"0152", x"0152", x"0152", x"0152", x"0152", x"0153", x"0153", x"0153", x"0153", x"0153", x"0153", x"0153", x"0153", x"0153", x"0153", x"0153", x"0153", x"0153", x"0154", x"0154", x"0154", x"0154", x"0154", x"0154", x"0154", x"0154", x"0154", x"0154", x"0154", x"0154", x"0154", x"0155", x"0155", x"0155", x"0155", x"0155", x"0155", x"0155", x"0155", x"0155", x"0155", x"0155", x"0155", x"0155", x"0155", x"0156", x"0156", x"0156", x"0156", x"0156", x"0156", x"0156", x"0156", x"0156", x"0156", x"0156", x"0156", x"0156", x"0157", x"0157", x"0157", x"0157", x"0157", x"0157", x"0157", x"0157", x"0157", x"0157", x"0157", x"0157", x"0157", x"0158", x"0158", x"0158", x"0158", x"0158", x"0158", x"0158", x"0158", x"0158", x"0158", x"0158", x"0158", x"0158", x"0159", x"0159", x"0159", x"0159", x"0159", x"0159", x"0159", x"0159", x"0159", x"0159", x"0159", x"0159", x"0159", x"015a", x"015a", x"015a", x"015a", x"015a", x"015a", x"015a", x"015a", x"015a", x"015a", x"015a", x"015a", x"015b", x"015b", x"015b", x"015b", x"015b", x"015b", x"015b", x"015b", x"015b", x"015b", x"015b", x"015b", x"015b", x"015c", x"015c", x"015c", x"015c", x"015c", x"015c", x"015c", x"015c", x"015c", x"015c", x"015c", x"015c", x"015c", x"015d", x"015d", x"015d", x"015d", x"015d", x"015d", x"015d", x"015d", x"015d", x"015d", x"015d", x"015d", x"015d", x"015e", x"015e", x"015e", x"015e", x"015e", x"015e", x"015e", x"015e", x"015e", x"015e", x"015e", x"015e", x"015e", x"015f", x"015f", x"015f", x"015f", x"015f", x"015f", x"015f", x"015f", x"015f", x"015f", x"015f", x"015f", x"015f", x"0160", x"0160", x"0160", x"0160", x"0160", x"0160", x"0160", x"0160", x"0160", x"0160", x"0160", x"0160", x"0161", x"0161", x"0161", x"0161", x"0161", x"0161", x"0161", x"0161", x"0161", x"0161", x"0161", x"0161", x"0161", x"0162", x"0162", x"0162", x"0162", x"0162", x"0162", x"0162", x"0162", x"0162", x"0162", x"0162", x"0162", x"0162", x"0163", x"0163", x"0163", x"0163", x"0163", x"0163", x"0163", x"0163", x"0163", x"0163", x"0163", x"0163", x"0164", x"0164", x"0164", x"0164", x"0164", x"0164", x"0164", x"0164", x"0164", x"0164", x"0164", x"0164", x"0164", x"0165", x"0165", x"0165", x"0165", x"0165", x"0165", x"0165", x"0165", x"0165", x"0165", x"0165", x"0165", x"0166", x"0166", x"0166", x"0166", x"0166", x"0166", x"0166", x"0166", x"0166", x"0166", x"0166", x"0166", x"0166", x"0167", x"0167", x"0167", x"0167", x"0167", x"0167", x"0167", x"0167", x"0167", x"0167", x"0167", x"0167", x"0168", x"0168", x"0168", x"0168", x"0168", x"0168", x"0168", x"0168", x"0168", x"0168", x"0168", x"0168", x"0168", x"0169", x"0169", x"0169", x"0169", x"0169", x"0169", x"0169", x"0169", x"0169", x"0169", x"0169", x"0169", x"016a", x"016a", x"016a", x"016a", x"016a", x"016a", x"016a", x"016a", x"016a", x"016a", x"016a", x"016a", x"016a", x"016b", x"016b", x"016b", x"016b", x"016b", x"016b", x"016b", x"016b", x"016b", x"016b", x"016b", x"016b", x"016c", x"016c", x"016c", x"016c", x"016c", x"016c", x"016c", x"016c", x"016c", x"016c", x"016c", x"016c", x"016d", x"016d", x"016d", x"016d", x"016d", x"016d", x"016d", x"016d", x"016d", x"016d", x"016d", x"016d", x"016d", x"016e", x"016e", x"016e", x"016e", x"016e", x"016e", x"016e", x"016e", x"016e", x"016e", x"016e", x"016e", x"016f", x"016f", x"016f", x"016f", x"016f", x"016f", x"016f", x"016f", x"016f", x"016f", x"016f", x"016f", x"0170", x"0170", x"0170", x"0170", x"0170", x"0170", x"0170", x"0170", x"0170", x"0170", x"0170", x"0170", x"0171", x"0171", x"0171", x"0171", x"0171", x"0171", x"0171", x"0171", x"0171", x"0171", x"0171", x"0171", x"0171", x"0172", x"0172", x"0172", x"0172", x"0172", x"0172", x"0172", x"0172", x"0172", x"0172", x"0172", x"0172", x"0173", x"0173", x"0173", x"0173", x"0173", x"0173", x"0173", x"0173", x"0173", x"0173", x"0173", x"0173", x"0174", x"0174", x"0174", x"0174", x"0174", x"0174", x"0174", x"0174", x"0174", x"0174", x"0174", x"0174", x"0175", x"0175", x"0175", x"0175", x"0175", x"0175", x"0175", x"0175", x"0175", x"0175", x"0175", x"0175", x"0176", x"0176", x"0176", x"0176", x"0176", x"0176", x"0176", x"0176", x"0176", x"0176", x"0176", x"0176", x"0177", x"0177", x"0177", x"0177", x"0177", x"0177", x"0177", x"0177", x"0177", x"0177", x"0177", x"0177", x"0178", x"0178", x"0178", x"0178", x"0178", x"0178", x"0178", x"0178", x"0178", x"0178", x"0178", x"0178", x"0179", x"0179", x"0179", x"0179", x"0179", x"0179", x"0179", x"0179", x"0179", x"0179", x"0179", x"0179", x"017a", x"017a", x"017a", x"017a", x"017a", x"017a", x"017a", x"017a", x"017a", x"017a", x"017a", x"017a", x"017b", x"017b", x"017b", x"017b", x"017b", x"017b", x"017b", x"017b", x"017b", x"017b", x"017b", x"017b", x"017c", x"017c", x"017c", x"017c", x"017c", x"017c", x"017c", x"017c", x"017c", x"017c", x"017c", x"017c", x"017d", x"017d", x"017d", x"017d", x"017d", x"017d", x"017d", x"017d", x"017d", x"017d", x"017d", x"017e", x"017e", x"017e", x"017e", x"017e", x"017e", x"017e", x"017e", x"017e", x"017e", x"017e", x"017e", x"017f", x"017f", x"017f", x"017f", x"017f", x"017f", x"017f", x"017f", x"017f", x"017f", x"017f", x"017f", x"0180", x"0180", x"0180", x"0180", x"0180", x"0180", x"0180", x"0180", x"0180", x"0180", x"0180", x"0180", x"0181", x"0181", x"0181", x"0181", x"0181", x"0181", x"0181", x"0181", x"0181", x"0181", x"0181", x"0181", x"0182", x"0182", x"0182", x"0182", x"0182", x"0182", x"0182", x"0182", x"0182", x"0182", x"0182", x"0183", x"0183", x"0183", x"0183", x"0183", x"0183", x"0183", x"0183", x"0183", x"0183", x"0183", x"0183", x"0184", x"0184", x"0184", x"0184", x"0184", x"0184", x"0184", x"0184", x"0184", x"0184", x"0184", x"0184", x"0185", x"0185", x"0185", x"0185", x"0185", x"0185", x"0185", x"0185", x"0185", x"0185", x"0185", x"0186", x"0186", x"0186", x"0186", x"0186", x"0186", x"0186", x"0186", x"0186", x"0186", x"0186", x"0186", x"0187", x"0187", x"0187", x"0187", x"0187", x"0187", x"0187", x"0187", x"0187", x"0187", x"0187", x"0188", x"0188", x"0188", x"0188", x"0188", x"0188", x"0188", x"0188", x"0188", x"0188", x"0188", x"0188", x"0189", x"0189", x"0189", x"0189", x"0189", x"0189", x"0189", x"0189", x"0189", x"0189", x"0189", x"018a", x"018a", x"018a", x"018a", x"018a", x"018a", x"018a", x"018a", x"018a", x"018a", x"018a", x"018a", x"018b", x"018b", x"018b", x"018b", x"018b", x"018b", x"018b", x"018b", x"018b", x"018b", x"018b", x"018c", x"018c", x"018c", x"018c", x"018c", x"018c", x"018c", x"018c", x"018c", x"018c", x"018c", x"018c", x"018d", x"018d", x"018d", x"018d", x"018d", x"018d", x"018d", x"018d", x"018d", x"018d", x"018d", x"018e", x"018e", x"018e", x"018e", x"018e", x"018e", x"018e", x"018e", x"018e", x"018e", x"018e", x"018e", x"018f", x"018f", x"018f", x"018f", x"018f", x"018f", x"018f", x"018f", x"018f", x"018f", x"018f", x"0190", x"0190", x"0190", x"0190", x"0190", x"0190", x"0190", x"0190", x"0190", x"0190", x"0190", x"0191", x"0191", x"0191", x"0191", x"0191", x"0191", x"0191", x"0191", x"0191", x"0191", x"0191", x"0191", x"0192", x"0192", x"0192", x"0192", x"0192", x"0192", x"0192", x"0192", x"0192", x"0192", x"0192", x"0193", x"0193", x"0193", x"0193", x"0193", x"0193", x"0193", x"0193", x"0193", x"0193", x"0193", x"0194", x"0194", x"0194", x"0194", x"0194", x"0194", x"0194", x"0194", x"0194", x"0194", x"0194", x"0195", x"0195", x"0195", x"0195", x"0195", x"0195", x"0195", x"0195", x"0195", x"0195", x"0195", x"0195", x"0196", x"0196", x"0196", x"0196", x"0196", x"0196", x"0196", x"0196", x"0196", x"0196", x"0196", x"0197", x"0197", x"0197", x"0197", x"0197", x"0197", x"0197", x"0197", x"0197", x"0197", x"0197", x"0198", x"0198", x"0198", x"0198", x"0198", x"0198", x"0198", x"0198", x"0198", x"0198", x"0198", x"0199", x"0199", x"0199", x"0199", x"0199", x"0199", x"0199", x"0199", x"0199", x"0199", x"0199", x"019a", x"019a", x"019a", x"019a", x"019a", x"019a", x"019a", x"019a", x"019a", x"019a", x"019a", x"019b", x"019b", x"019b", x"019b", x"019b", x"019b", x"019b", x"019b", x"019b", x"019b", x"019b", x"019c", x"019c", x"019c", x"019c", x"019c", x"019c", x"019c", x"019c", x"019c", x"019c", x"019c", x"019d", x"019d", x"019d", x"019d", x"019d", x"019d", x"019d", x"019d", x"019d", x"019d", x"019d", x"019e", x"019e", x"019e", x"019e", x"019e", x"019e", x"019e", x"019e", x"019e", x"019e", x"019e", x"019f", x"019f", x"019f", x"019f", x"019f", x"019f", x"019f", x"019f", x"019f", x"019f", x"019f", x"01a0", x"01a0", x"01a0", x"01a0", x"01a0", x"01a0", x"01a0", x"01a0", x"01a0", x"01a0", x"01a0", x"01a1", x"01a1", x"01a1", x"01a1", x"01a1", x"01a1", x"01a1", x"01a1", x"01a1", x"01a1", x"01a1", x"01a2", x"01a2", x"01a2", x"01a2", x"01a2", x"01a2", x"01a2", x"01a2", x"01a2", x"01a2", x"01a2", x"01a3", x"01a3", x"01a3", x"01a3", x"01a3", x"01a3", x"01a3", x"01a3", x"01a3", x"01a3", x"01a3", x"01a4", x"01a4", x"01a4", x"01a4", x"01a4", x"01a4", x"01a4", x"01a4", x"01a4", x"01a4", x"01a4", x"01a5", x"01a5", x"01a5", x"01a5", x"01a5", x"01a5", x"01a5", x"01a5", x"01a5", x"01a5", x"01a5", x"01a6", x"01a6", x"01a6", x"01a6", x"01a6", x"01a6", x"01a6", x"01a6", x"01a6", x"01a6", x"01a6", x"01a7", x"01a7", x"01a7", x"01a7", x"01a7", x"01a7", x"01a7", x"01a7", x"01a7", x"01a7", x"01a8", x"01a8", x"01a8", x"01a8", x"01a8", x"01a8", x"01a8", x"01a8", x"01a8", x"01a8", x"01a8", x"01a9", x"01a9", x"01a9", x"01a9", x"01a9", x"01a9", x"01a9", x"01a9", x"01a9", x"01a9", x"01a9", x"01aa", x"01aa", x"01aa", x"01aa", x"01aa", x"01aa", x"01aa", x"01aa", x"01aa", x"01aa", x"01aa", x"01ab", x"01ab", x"01ab", x"01ab", x"01ab", x"01ab", x"01ab", x"01ab", x"01ab", x"01ab", x"01ac", x"01ac", x"01ac", x"01ac", x"01ac", x"01ac", x"01ac", x"01ac", x"01ac", x"01ac", x"01ac", x"01ad", x"01ad", x"01ad", x"01ad", x"01ad", x"01ad", x"01ad", x"01ad", x"01ad", x"01ad", x"01ad", x"01ae", x"01ae", x"01ae", x"01ae", x"01ae", x"01ae", x"01ae", x"01ae", x"01ae", x"01ae", x"01af", x"01af", x"01af", x"01af", x"01af", x"01af", x"01af", x"01af", x"01af", x"01af", x"01af", x"01b0", x"01b0", x"01b0", x"01b0", x"01b0", x"01b0", x"01b0", x"01b0", x"01b0", x"01b0", x"01b1", x"01b1", x"01b1", x"01b1", x"01b1", x"01b1", x"01b1", x"01b1", x"01b1", x"01b1", x"01b1", x"01b2", x"01b2", x"01b2", x"01b2", x"01b2", x"01b2", x"01b2", x"01b2", x"01b2", x"01b2", x"01b2", x"01b3", x"01b3", x"01b3", x"01b3", x"01b3", x"01b3", x"01b3", x"01b3", x"01b3", x"01b3", x"01b4", x"01b4", x"01b4", x"01b4", x"01b4", x"01b4", x"01b4", x"01b4", x"01b4", x"01b4", x"01b4", x"01b5", x"01b5", x"01b5", x"01b5", x"01b5", x"01b5", x"01b5", x"01b5", x"01b5", x"01b5", x"01b6", x"01b6", x"01b6", x"01b6", x"01b6", x"01b6", x"01b6", x"01b6", x"01b6", x"01b6", x"01b6", x"01b7", x"01b7", x"01b7", x"01b7", x"01b7", x"01b7", x"01b7", x"01b7", x"01b7", x"01b7", x"01b8", x"01b8", x"01b8", x"01b8", x"01b8", x"01b8", x"01b8", x"01b8", x"01b8", x"01b8", x"01b9", x"01b9", x"01b9", x"01b9", x"01b9", x"01b9", x"01b9", x"01b9", x"01b9", x"01b9", x"01b9", x"01ba", x"01ba", x"01ba", x"01ba", x"01ba", x"01ba", x"01ba", x"01ba", x"01ba", x"01ba", x"01bb", x"01bb", x"01bb", x"01bb", x"01bb", x"01bb", x"01bb", x"01bb", x"01bb", x"01bb", x"01bb", x"01bc", x"01bc", x"01bc", x"01bc", x"01bc", x"01bc", x"01bc", x"01bc", x"01bc", x"01bc", x"01bd", x"01bd", x"01bd", x"01bd", x"01bd", x"01bd", x"01bd", x"01bd", x"01bd", x"01bd", x"01be", x"01be", x"01be", x"01be", x"01be", x"01be", x"01be", x"01be", x"01be", x"01be", x"01bf", x"01bf", x"01bf", x"01bf", x"01bf", x"01bf", x"01bf", x"01bf", x"01bf", x"01bf", x"01bf", x"01c0", x"01c0", x"01c0", x"01c0", x"01c0", x"01c0", x"01c0", x"01c0", x"01c0", x"01c0", x"01c1", x"01c1", x"01c1", x"01c1", x"01c1", x"01c1", x"01c1", x"01c1", x"01c1", x"01c1", x"01c2", x"01c2", x"01c2", x"01c2", x"01c2", x"01c2", x"01c2", x"01c2", x"01c2", x"01c2", x"01c3", x"01c3", x"01c3", x"01c3", x"01c3", x"01c3", x"01c3", x"01c3", x"01c3", x"01c3", x"01c3", x"01c4", x"01c4", x"01c4", x"01c4", x"01c4", x"01c4", x"01c4", x"01c4", x"01c4", x"01c4", x"01c5", x"01c5", x"01c5", x"01c5", x"01c5", x"01c5", x"01c5", x"01c5", x"01c5", x"01c5", x"01c6", x"01c6", x"01c6", x"01c6", x"01c6", x"01c6", x"01c6", x"01c6", x"01c6", x"01c6", x"01c7", x"01c7", x"01c7", x"01c7", x"01c7", x"01c7", x"01c7", x"01c7", x"01c7", x"01c7", x"01c8", x"01c8", x"01c8", x"01c8", x"01c8", x"01c8", x"01c8", x"01c8", x"01c8", x"01c8", x"01c9", x"01c9", x"01c9", x"01c9", x"01c9", x"01c9", x"01c9", x"01c9", x"01c9", x"01c9", x"01ca", x"01ca", x"01ca", x"01ca", x"01ca", x"01ca", x"01ca", x"01ca", x"01ca", x"01ca", x"01cb", x"01cb", x"01cb", x"01cb", x"01cb", x"01cb", x"01cb", x"01cb", x"01cb", x"01cb", x"01cb", x"01cc", x"01cc", x"01cc", x"01cc", x"01cc", x"01cc", x"01cc", x"01cc", x"01cc", x"01cc", x"01cd", x"01cd", x"01cd", x"01cd", x"01cd", x"01cd", x"01cd", x"01cd", x"01cd", x"01cd", x"01ce", x"01ce", x"01ce", x"01ce", x"01ce", x"01ce", x"01ce", x"01ce", x"01ce", x"01ce", x"01cf", x"01cf", x"01cf", x"01cf", x"01cf", x"01cf", x"01cf", x"01cf", x"01cf", x"01d0", x"01d0", x"01d0", x"01d0", x"01d0", x"01d0", x"01d0", x"01d0", x"01d0", x"01d0", x"01d1", x"01d1", x"01d1", x"01d1", x"01d1", x"01d1", x"01d1", x"01d1", x"01d1", x"01d1", x"01d2", x"01d2", x"01d2", x"01d2", x"01d2", x"01d2", x"01d2", x"01d2", x"01d2", x"01d2", x"01d3", x"01d3", x"01d3", x"01d3", x"01d3", x"01d3", x"01d3", x"01d3", x"01d3", x"01d3", x"01d4", x"01d4", x"01d4", x"01d4", x"01d4", x"01d4", x"01d4", x"01d4", x"01d4", x"01d4", x"01d5", x"01d5", x"01d5", x"01d5", x"01d5", x"01d5", x"01d5", x"01d5", x"01d5", x"01d5", x"01d6", x"01d6", x"01d6", x"01d6", x"01d6", x"01d6", x"01d6", x"01d6", x"01d6", x"01d6", x"01d7", x"01d7", x"01d7", x"01d7", x"01d7", x"01d7", x"01d7", x"01d7", x"01d7", x"01d7", x"01d8", x"01d8", x"01d8", x"01d8", x"01d8", x"01d8", x"01d8", x"01d8", x"01d8", x"01d9", x"01d9", x"01d9", x"01d9", x"01d9", x"01d9", x"01d9", x"01d9", x"01d9", x"01d9", x"01da", x"01da", x"01da", x"01da", x"01da", x"01da", x"01da", x"01da", x"01da", x"01da", x"01db", x"01db", x"01db", x"01db", x"01db", x"01db", x"01db", x"01db", x"01db", x"01db", x"01dc", x"01dc", x"01dc", x"01dc", x"01dc", x"01dc", x"01dc", x"01dc", x"01dc", x"01dd", x"01dd", x"01dd", x"01dd", x"01dd", x"01dd", x"01dd", x"01dd", x"01dd", x"01dd", x"01de", x"01de", x"01de", x"01de", x"01de", x"01de", x"01de", x"01de", x"01de", x"01de", x"01df", x"01df", x"01df", x"01df", x"01df", x"01df", x"01df", x"01df", x"01df", x"01e0", x"01e0", x"01e0", x"01e0", x"01e0", x"01e0", x"01e0", x"01e0", x"01e0", x"01e0", x"01e1", x"01e1", x"01e1", x"01e1", x"01e1", x"01e1", x"01e1", x"01e1", x"01e1", x"01e1", x"01e2", x"01e2", x"01e2", x"01e2", x"01e2", x"01e2", x"01e2", x"01e2", x"01e2", x"01e3", x"01e3", x"01e3", x"01e3", x"01e3", x"01e3", x"01e3", x"01e3", x"01e3", x"01e3", x"01e4", x"01e4", x"01e4", x"01e4", x"01e4", x"01e4", x"01e4", x"01e4", x"01e4", x"01e4", x"01e5", x"01e5", x"01e5", x"01e5", x"01e5", x"01e5", x"01e5", x"01e5", x"01e5", x"01e6", x"01e6", x"01e6", x"01e6", x"01e6", x"01e6", x"01e6", x"01e6", x"01e6", x"01e6", x"01e7", x"01e7", x"01e7", x"01e7", x"01e7", x"01e7", x"01e7", x"01e7", x"01e7", x"01e8", x"01e8", x"01e8", x"01e8", x"01e8", x"01e8", x"01e8", x"01e8", x"01e8", x"01e8", x"01e9", x"01e9", x"01e9", x"01e9", x"01e9", x"01e9", x"01e9", x"01e9", x"01e9", x"01ea", x"01ea", x"01ea", x"01ea", x"01ea", x"01ea", x"01ea", x"01ea", x"01ea", x"01ea", x"01eb", x"01eb", x"01eb", x"01eb", x"01eb", x"01eb", x"01eb", x"01eb", x"01eb", x"01ec", x"01ec", x"01ec", x"01ec", x"01ec", x"01ec", x"01ec", x"01ec", x"01ec", x"01ec", x"01ed", x"01ed", x"01ed", x"01ed", x"01ed", x"01ed", x"01ed", x"01ed", x"01ed", x"01ee", x"01ee", x"01ee", x"01ee", x"01ee", x"01ee", x"01ee", x"01ee", x"01ee", x"01ef", x"01ef", x"01ef", x"01ef", x"01ef", x"01ef", x"01ef", x"01ef", x"01ef", x"01ef", x"01f0", x"01f0", x"01f0", x"01f0", x"01f0", x"01f0", x"01f0", x"01f0", x"01f0", x"01f1", x"01f1", x"01f1", x"01f1", x"01f1", x"01f1", x"01f1", x"01f1", x"01f1", x"01f1", x"01f2", x"01f2", x"01f2", x"01f2", x"01f2", x"01f2", x"01f2", x"01f2", x"01f2", x"01f3", x"01f3", x"01f3", x"01f3", x"01f3", x"01f3", x"01f3", x"01f3", x"01f3", x"01f4", x"01f4", x"01f4", x"01f4", x"01f4", x"01f4", x"01f4", x"01f4", x"01f4", x"01f4", x"01f5", x"01f5", x"01f5", x"01f5", x"01f5", x"01f5", x"01f5", x"01f5", x"01f5", x"01f6", x"01f6", x"01f6", x"01f6", x"01f6", x"01f6", x"01f6", x"01f6", x"01f6", x"01f7", x"01f7", x"01f7", x"01f7", x"01f7", x"01f7", x"01f7", x"01f7", x"01f7", x"01f7", x"01f8", x"01f8", x"01f8", x"01f8", x"01f8", x"01f8", x"01f8", x"01f8", x"01f8", x"01f9", x"01f9", x"01f9", x"01f9", x"01f9", x"01f9", x"01f9", x"01f9", x"01f9", x"01fa", x"01fa", x"01fa", x"01fa", x"01fa", x"01fa", x"01fa", x"01fa", x"01fa", x"01fb", x"01fb", x"01fb", x"01fb", x"01fb", x"01fb", x"01fb", x"01fb", x"01fb", x"01fc", x"01fc", x"01fc", x"01fc", x"01fc", x"01fc", x"01fc", x"01fc", x"01fc", x"01fc", x"01fd", x"01fd", x"01fd", x"01fd", x"01fd", x"01fd", x"01fd", x"01fd", x"01fd", x"01fe", x"01fe", x"01fe", x"01fe", x"01fe", x"01fe", x"01fe", x"01fe", x"01fe", x"01ff", x"01ff", x"01ff", x"01ff", x"01ff", x"01ff", x"01ff", x"01ff", x"01ff", x"0200", x"0200", x"0200", x"0200", x"0200", x"0200", x"0200", x"0200", x"0200", x"0201", x"0201", x"0201", x"0201", x"0201", x"0201", x"0201", x"0201", x"0201", x"0202", x"0202", x"0202", x"0202", x"0202", x"0202", x"0202", x"0202", x"0202", x"0202", x"0203", x"0203", x"0203", x"0203", x"0203", x"0203", x"0203", x"0203", x"0203", x"0204", x"0204", x"0204", x"0204", x"0204", x"0204", x"0204", x"0204", x"0204", x"0205", x"0205", x"0205", x"0205", x"0205", x"0205", x"0205", x"0205", x"0205", x"0206", x"0206", x"0206", x"0206", x"0206", x"0206", x"0206", x"0206", x"0206", x"0207", x"0207", x"0207", x"0207", x"0207", x"0207", x"0207", x"0207", x"0207", x"0208", x"0208", x"0208", x"0208", x"0208", x"0208", x"0208", x"0208", x"0208", x"0209", x"0209", x"0209", x"0209", x"0209", x"0209", x"0209", x"0209", x"0209", x"020a", x"020a", x"020a", x"020a", x"020a", x"020a", x"020a", x"020a", x"020a", x"020b", x"020b", x"020b", x"020b", x"020b", x"020b", x"020b", x"020b", x"020b", x"020c", x"020c", x"020c", x"020c", x"020c", x"020c", x"020c", x"020c", x"020c", x"020d", x"020d", x"020d", x"020d", x"020d", x"020d", x"020d", x"020d", x"020d", x"020e", x"020e", x"020e", x"020e", x"020e", x"020e", x"020e", x"020e", x"020e", x"020f", x"020f", x"020f", x"020f", x"020f", x"020f", x"020f", x"020f", x"020f", x"0210", x"0210", x"0210", x"0210", x"0210", x"0210", x"0210", x"0210", x"0211", x"0211", x"0211", x"0211", x"0211", x"0211", x"0211", x"0211", x"0211", x"0212", x"0212", x"0212", x"0212", x"0212", x"0212", x"0212", x"0212", x"0212", x"0213", x"0213", x"0213", x"0213", x"0213", x"0213", x"0213", x"0213", x"0213", x"0214", x"0214", x"0214", x"0214", x"0214", x"0214", x"0214", x"0214", x"0214", x"0215", x"0215", x"0215", x"0215", x"0215", x"0215", x"0215", x"0215", x"0215", x"0216", x"0216", x"0216", x"0216", x"0216", x"0216", x"0216", x"0216", x"0216", x"0217", x"0217", x"0217", x"0217", x"0217", x"0217", x"0217", x"0217", x"0218", x"0218", x"0218", x"0218", x"0218", x"0218", x"0218", x"0218", x"0218", x"0219", x"0219", x"0219", x"0219", x"0219", x"0219", x"0219", x"0219", x"0219", x"021a", x"021a", x"021a", x"021a", x"021a", x"021a", x"021a", x"021a", x"021a", x"021b", x"021b", x"021b", x"021b", x"021b", x"021b", x"021b", x"021b", x"021c", x"021c", x"021c", x"021c", x"021c", x"021c", x"021c", x"021c", x"021c", x"021d", x"021d", x"021d", x"021d", x"021d", x"021d", x"021d", x"021d", x"021d", x"021e", x"021e", x"021e", x"021e", x"021e", x"021e", x"021e", x"021e", x"021e", x"021f", x"021f", x"021f", x"021f", x"021f", x"021f", x"021f", x"021f", x"0220", x"0220", x"0220", x"0220", x"0220", x"0220", x"0220", x"0220", x"0220", x"0221", x"0221", x"0221", x"0221", x"0221", x"0221", x"0221", x"0221", x"0221", x"0222", x"0222", x"0222", x"0222", x"0222", x"0222", x"0222", x"0222", x"0223", x"0223", x"0223", x"0223", x"0223", x"0223", x"0223", x"0223", x"0223", x"0224", x"0224", x"0224", x"0224", x"0224", x"0224", x"0224", x"0224", x"0224", x"0225", x"0225", x"0225", x"0225", x"0225", x"0225", x"0225", x"0225", x"0226", x"0226", x"0226", x"0226", x"0226", x"0226", x"0226", x"0226", x"0226", x"0227", x"0227", x"0227", x"0227", x"0227", x"0227", x"0227", x"0227", x"0228", x"0228", x"0228", x"0228", x"0228", x"0228", x"0228", x"0228", x"0228", x"0229", x"0229", x"0229", x"0229", x"0229", x"0229", x"0229", x"0229", x"022a", x"022a", x"022a", x"022a", x"022a", x"022a", x"022a", x"022a", x"022a", x"022b", x"022b", x"022b", x"022b", x"022b", x"022b", x"022b", x"022b", x"022c", x"022c", x"022c", x"022c", x"022c", x"022c", x"022c", x"022c", x"022c", x"022d", x"022d", x"022d", x"022d", x"022d", x"022d", x"022d", x"022d", x"022d", x"022e", x"022e", x"022e", x"022e", x"022e", x"022e", x"022e", x"022e", x"022f", x"022f", x"022f", x"022f", x"022f", x"022f", x"022f", x"022f", x"0230", x"0230", x"0230", x"0230", x"0230", x"0230", x"0230", x"0230", x"0230", x"0231", x"0231", x"0231", x"0231", x"0231", x"0231", x"0231", x"0231", x"0232", x"0232", x"0232", x"0232", x"0232", x"0232", x"0232", x"0232", x"0232", x"0233", x"0233", x"0233", x"0233", x"0233", x"0233", x"0233", x"0233", x"0234", x"0234", x"0234", x"0234", x"0234", x"0234", x"0234", x"0234", x"0234", x"0235", x"0235", x"0235", x"0235", x"0235", x"0235", x"0235", x"0235", x"0236", x"0236", x"0236", x"0236", x"0236", x"0236", x"0236", x"0236", x"0237", x"0237", x"0237", x"0237", x"0237", x"0237", x"0237", x"0237", x"0237", x"0238", x"0238", x"0238", x"0238", x"0238", x"0238", x"0238", x"0238", x"0239", x"0239", x"0239", x"0239", x"0239", x"0239", x"0239", x"0239", x"0239", x"023a", x"023a", x"023a", x"023a", x"023a", x"023a", x"023a", x"023a", x"023b", x"023b", x"023b", x"023b", x"023b", x"023b", x"023b", x"023b", x"023c", x"023c", x"023c", x"023c", x"023c", x"023c", x"023c", x"023c", x"023c", x"023d", x"023d", x"023d", x"023d", x"023d", x"023d", x"023d", x"023d", x"023e", x"023e", x"023e", x"023e", x"023e", x"023e", x"023e", x"023e", x"023f", x"023f", x"023f", x"023f", x"023f", x"023f", x"023f", x"023f", x"0240", x"0240", x"0240", x"0240", x"0240", x"0240", x"0240", x"0240", x"0240", x"0241", x"0241", x"0241", x"0241", x"0241", x"0241", x"0241", x"0241", x"0242", x"0242", x"0242", x"0242", x"0242", x"0242", x"0242", x"0242", x"0243", x"0243", x"0243", x"0243", x"0243", x"0243", x"0243", x"0243", x"0244", x"0244", x"0244", x"0244", x"0244", x"0244", x"0244", x"0244", x"0244", x"0245", x"0245", x"0245", x"0245", x"0245", x"0245", x"0245", x"0245", x"0246", x"0246", x"0246", x"0246", x"0246", x"0246", x"0246", x"0246", x"0247", x"0247", x"0247", x"0247", x"0247", x"0247", x"0247", x"0247", x"0248", x"0248", x"0248", x"0248", x"0248", x"0248", x"0248", x"0248", x"0249", x"0249", x"0249", x"0249", x"0249", x"0249", x"0249", x"0249", x"0249", x"024a", x"024a", x"024a", x"024a", x"024a", x"024a", x"024a", x"024a", x"024b", x"024b", x"024b", x"024b", x"024b", x"024b", x"024b", x"024b", x"024c", x"024c", x"024c", x"024c", x"024c", x"024c", x"024c", x"024c", x"024d", x"024d", x"024d", x"024d", x"024d", x"024d", x"024d", x"024d", x"024e", x"024e", x"024e", x"024e", x"024e", x"024e", x"024e", x"024e", x"024f", x"024f", x"024f", x"024f", x"024f", x"024f", x"024f", x"024f", x"0250", x"0250", x"0250", x"0250", x"0250", x"0250", x"0250", x"0250", x"0251", x"0251", x"0251", x"0251", x"0251", x"0251", x"0251", x"0251", x"0251", x"0252", x"0252", x"0252", x"0252", x"0252", x"0252", x"0252", x"0252", x"0253", x"0253", x"0253", x"0253", x"0253", x"0253", x"0253", x"0253", x"0254", x"0254", x"0254", x"0254", x"0254", x"0254", x"0254", x"0254", x"0255", x"0255", x"0255", x"0255", x"0255", x"0255", x"0255", x"0255", x"0256", x"0256", x"0256", x"0256", x"0256", x"0256", x"0256", x"0256", x"0257", x"0257", x"0257", x"0257", x"0257", x"0257", x"0257", x"0257", x"0258", x"0258", x"0258", x"0258", x"0258", x"0258", x"0258", x"0258", x"0259", x"0259", x"0259", x"0259", x"0259", x"0259", x"0259", x"0259", x"025a", x"025a", x"025a", x"025a", x"025a", x"025a", x"025a", x"025a", x"025b", x"025b", x"025b", x"025b", x"025b", x"025b", x"025b", x"025b", x"025c", x"025c", x"025c", x"025c", x"025c", x"025c", x"025c", x"025c", x"025d", x"025d", x"025d", x"025d", x"025d", x"025d", x"025d", x"025e", x"025e", x"025e", x"025e", x"025e", x"025e", x"025e", x"025e", x"025f", x"025f", x"025f", x"025f", x"025f", x"025f", x"025f", x"025f", x"0260", x"0260", x"0260", x"0260", x"0260", x"0260", x"0260", x"0260", x"0261", x"0261", x"0261", x"0261", x"0261", x"0261", x"0261", x"0261", x"0262", x"0262", x"0262", x"0262", x"0262", x"0262", x"0262", x"0262", x"0263", x"0263", x"0263", x"0263", x"0263", x"0263", x"0263", x"0263", x"0264", x"0264", x"0264", x"0264", x"0264", x"0264", x"0264", x"0264", x"0265", x"0265", x"0265", x"0265", x"0265", x"0265", x"0265", x"0265", x"0266", x"0266", x"0266", x"0266", x"0266", x"0266", x"0266", x"0267", x"0267", x"0267", x"0267", x"0267", x"0267", x"0267", x"0267", x"0268", x"0268", x"0268", x"0268", x"0268", x"0268", x"0268", x"0268", x"0269", x"0269", x"0269", x"0269", x"0269", x"0269", x"0269", x"0269", x"026a", x"026a", x"026a", x"026a", x"026a", x"026a", x"026a", x"026a", x"026b", x"026b", x"026b", x"026b", x"026b", x"026b", x"026b", x"026b", x"026c", x"026c", x"026c", x"026c", x"026c", x"026c", x"026c", x"026d", x"026d", x"026d", x"026d", x"026d", x"026d", x"026d", x"026d", x"026e", x"026e", x"026e", x"026e", x"026e", x"026e", x"026e", x"026e", x"026f", x"026f", x"026f", x"026f", x"026f", x"026f", x"026f", x"026f", x"0270", x"0270", x"0270", x"0270", x"0270", x"0270", x"0270", x"0271", x"0271", x"0271", x"0271", x"0271", x"0271", x"0271", x"0271", x"0272", x"0272", x"0272", x"0272", x"0272", x"0272", x"0272", x"0272", x"0273", x"0273", x"0273", x"0273", x"0273", x"0273", x"0273", x"0274", x"0274", x"0274", x"0274", x"0274", x"0274", x"0274", x"0274", x"0275", x"0275", x"0275", x"0275", x"0275", x"0275", x"0275", x"0275", x"0276", x"0276", x"0276", x"0276", x"0276", x"0276", x"0276", x"0276", x"0277", x"0277", x"0277", x"0277", x"0277", x"0277", x"0277", x"0278", x"0278", x"0278", x"0278", x"0278", x"0278", x"0278", x"0278", x"0279", x"0279", x"0279", x"0279", x"0279", x"0279", x"0279", x"0279", x"027a", x"027a", x"027a", x"027a", x"027a", x"027a", x"027a", x"027b", x"027b", x"027b", x"027b", x"027b", x"027b", x"027b", x"027b", x"027c", x"027c", x"027c", x"027c", x"027c", x"027c", x"027c", x"027d", x"027d", x"027d", x"027d", x"027d", x"027d", x"027d", x"027d", x"027e", x"027e", x"027e", x"027e", x"027e", x"027e", x"027e", x"027e", x"027f", x"027f", x"027f", x"027f", x"027f", x"027f", x"027f", x"0280", x"0280", x"0280", x"0280", x"0280", x"0280", x"0280", x"0280", x"0281", x"0281", x"0281", x"0281", x"0281", x"0281", x"0281", x"0282", x"0282", x"0282", x"0282", x"0282", x"0282", x"0282", x"0282", x"0283", x"0283", x"0283", x"0283", x"0283", x"0283", x"0283", x"0284", x"0284", x"0284", x"0284", x"0284", x"0284", x"0284", x"0284", x"0285", x"0285", x"0285", x"0285", x"0285", x"0285", x"0285", x"0285", x"0286", x"0286", x"0286", x"0286", x"0286", x"0286", x"0286", x"0287", x"0287", x"0287", x"0287", x"0287", x"0287", x"0287", x"0287", x"0288", x"0288", x"0288", x"0288", x"0288", x"0288", x"0288", x"0289", x"0289", x"0289", x"0289", x"0289", x"0289", x"0289", x"0289", x"028a", x"028a", x"028a", x"028a", x"028a", x"028a", x"028a", x"028b", x"028b", x"028b", x"028b", x"028b", x"028b", x"028b", x"028b", x"028c", x"028c", x"028c", x"028c", x"028c", x"028c", x"028c", x"028d", x"028d", x"028d", x"028d", x"028d", x"028d", x"028d", x"028e", x"028e", x"028e", x"028e", x"028e", x"028e", x"028e", x"028e", x"028f", x"028f", x"028f", x"028f", x"028f", x"028f", x"028f", x"0290", x"0290", x"0290", x"0290", x"0290", x"0290", x"0290", x"0290", x"0291", x"0291", x"0291", x"0291", x"0291", x"0291", x"0291", x"0292", x"0292", x"0292", x"0292", x"0292", x"0292", x"0292", x"0292", x"0293", x"0293", x"0293", x"0293", x"0293", x"0293", x"0293", x"0294", x"0294", x"0294", x"0294", x"0294", x"0294", x"0294", x"0295", x"0295", x"0295", x"0295", x"0295", x"0295", x"0295", x"0295", x"0296", x"0296", x"0296", x"0296", x"0296", x"0296", x"0296", x"0297", x"0297", x"0297", x"0297", x"0297", x"0297", x"0297", x"0297", x"0298", x"0298", x"0298", x"0298", x"0298", x"0298", x"0298", x"0299", x"0299", x"0299", x"0299", x"0299", x"0299", x"0299", x"029a", x"029a", x"029a", x"029a", x"029a", x"029a", x"029a", x"029a", x"029b", x"029b", x"029b", x"029b", x"029b", x"029b", x"029b", x"029c", x"029c", x"029c", x"029c", x"029c", x"029c", x"029c", x"029d", x"029d", x"029d", x"029d", x"029d", x"029d", x"029d", x"029d", x"029e", x"029e", x"029e", x"029e", x"029e", x"029e", x"029e", x"029f", x"029f", x"029f", x"029f", x"029f", x"029f", x"029f", x"02a0", x"02a0", x"02a0", x"02a0", x"02a0", x"02a0", x"02a0", x"02a1", x"02a1", x"02a1", x"02a1", x"02a1", x"02a1", x"02a1", x"02a1", x"02a2", x"02a2", x"02a2", x"02a2", x"02a2", x"02a2", x"02a2", x"02a3", x"02a3", x"02a3", x"02a3", x"02a3", x"02a3", x"02a3", x"02a4", x"02a4", x"02a4", x"02a4", x"02a4", x"02a4", x"02a4", x"02a4", x"02a5", x"02a5", x"02a5", x"02a5", x"02a5", x"02a5", x"02a5", x"02a6", x"02a6", x"02a6", x"02a6", x"02a6", x"02a6", x"02a6", x"02a7", x"02a7", x"02a7", x"02a7", x"02a7", x"02a7", x"02a7", x"02a8", x"02a8", x"02a8", x"02a8", x"02a8", x"02a8", x"02a8", x"02a9", x"02a9", x"02a9", x"02a9", x"02a9", x"02a9", x"02a9", x"02a9", x"02aa", x"02aa", x"02aa", x"02aa", x"02aa", x"02aa", x"02aa", x"02ab", x"02ab", x"02ab", x"02ab", x"02ab", x"02ab", x"02ab", x"02ac", x"02ac", x"02ac", x"02ac", x"02ac", x"02ac", x"02ac", x"02ad", x"02ad", x"02ad", x"02ad", x"02ad", x"02ad", x"02ad", x"02ae", x"02ae", x"02ae", x"02ae", x"02ae", x"02ae", x"02ae", x"02ae", x"02af", x"02af", x"02af", x"02af", x"02af", x"02af", x"02af", x"02b0", x"02b0", x"02b0", x"02b0", x"02b0", x"02b0", x"02b0", x"02b1", x"02b1", x"02b1", x"02b1", x"02b1", x"02b1", x"02b1", x"02b2", x"02b2", x"02b2", x"02b2", x"02b2", x"02b2", x"02b2", x"02b3", x"02b3", x"02b3", x"02b3", x"02b3", x"02b3", x"02b3", x"02b4", x"02b4", x"02b4", x"02b4", x"02b4", x"02b4", x"02b4", x"02b5", x"02b5", x"02b5", x"02b5", x"02b5", x"02b5", x"02b5", x"02b5", x"02b6", x"02b6", x"02b6", x"02b6", x"02b6", x"02b6", x"02b6", x"02b7", x"02b7", x"02b7", x"02b7", x"02b7", x"02b7", x"02b7", x"02b8", x"02b8", x"02b8", x"02b8", x"02b8", x"02b8", x"02b8", x"02b9", x"02b9", x"02b9", x"02b9", x"02b9", x"02b9", x"02b9", x"02ba", x"02ba", x"02ba", x"02ba", x"02ba", x"02ba", x"02ba", x"02bb", x"02bb", x"02bb", x"02bb", x"02bb", x"02bb", x"02bb", x"02bc", x"02bc", x"02bc", x"02bc", x"02bc", x"02bc", x"02bc", x"02bd", x"02bd", x"02bd", x"02bd", x"02bd", x"02bd", x"02bd", x"02be", x"02be", x"02be", x"02be", x"02be", x"02be", x"02be", x"02bf", x"02bf", x"02bf", x"02bf", x"02bf", x"02bf", x"02bf", x"02c0", x"02c0", x"02c0", x"02c0", x"02c0", x"02c0", x"02c0", x"02c1", x"02c1", x"02c1", x"02c1", x"02c1", x"02c1", x"02c1", x"02c2", x"02c2", x"02c2", x"02c2", x"02c2", x"02c2", x"02c2", x"02c3", x"02c3", x"02c3", x"02c3", x"02c3", x"02c3", x"02c3", x"02c4", x"02c4", x"02c4", x"02c4", x"02c4", x"02c4", x"02c4", x"02c5", x"02c5", x"02c5", x"02c5", x"02c5", x"02c5", x"02c5", x"02c6", x"02c6", x"02c6", x"02c6", x"02c6", x"02c6", x"02c6", x"02c7", x"02c7", x"02c7", x"02c7", x"02c7", x"02c7", x"02c7", x"02c8", x"02c8", x"02c8", x"02c8", x"02c8", x"02c8", x"02c8", x"02c9", x"02c9", x"02c9", x"02c9", x"02c9", x"02c9", x"02c9", x"02ca", x"02ca", x"02ca", x"02ca", x"02ca", x"02ca", x"02ca", x"02cb", x"02cb", x"02cb", x"02cb", x"02cb", x"02cb", x"02cb", x"02cc", x"02cc", x"02cc", x"02cc", x"02cc", x"02cc", x"02cc", x"02cd", x"02cd", x"02cd", x"02cd", x"02cd", x"02cd", x"02cd", x"02ce", x"02ce", x"02ce", x"02ce", x"02ce", x"02ce", x"02ce", x"02cf", x"02cf", x"02cf", x"02cf", x"02cf", x"02cf", x"02cf", x"02d0", x"02d0", x"02d0", x"02d0", x"02d0", x"02d0", x"02d1", x"02d1", x"02d1", x"02d1", x"02d1", x"02d1", x"02d1", x"02d2", x"02d2", x"02d2", x"02d2", x"02d2", x"02d2", x"02d2", x"02d3", x"02d3", x"02d3", x"02d3", x"02d3", x"02d3", x"02d3", x"02d4", x"02d4", x"02d4", x"02d4", x"02d4", x"02d4", x"02d4", x"02d5", x"02d5", x"02d5", x"02d5", x"02d5", x"02d5", x"02d5", x"02d6", x"02d6", x"02d6", x"02d6", x"02d6", x"02d6", x"02d6", x"02d7", x"02d7", x"02d7", x"02d7", x"02d7", x"02d7", x"02d7", x"02d8", x"02d8", x"02d8", x"02d8", x"02d8", x"02d8", x"02d9", x"02d9", x"02d9", x"02d9", x"02d9", x"02d9", x"02d9", x"02da", x"02da", x"02da", x"02da", x"02da", x"02da", x"02da", x"02db", x"02db", x"02db", x"02db", x"02db", x"02db", x"02db", x"02dc", x"02dc", x"02dc", x"02dc", x"02dc", x"02dc", x"02dc", x"02dd", x"02dd", x"02dd", x"02dd", x"02dd", x"02dd", x"02de", x"02de", x"02de", x"02de", x"02de", x"02de", x"02de", x"02df", x"02df", x"02df", x"02df", x"02df", x"02df", x"02df", x"02e0", x"02e0", x"02e0", x"02e0", x"02e0", x"02e0", x"02e0", x"02e1", x"02e1", x"02e1", x"02e1", x"02e1", x"02e1", x"02e1", x"02e2", x"02e2", x"02e2", x"02e2", x"02e2", x"02e2", x"02e3", x"02e3", x"02e3", x"02e3", x"02e3", x"02e3", x"02e3", x"02e4", x"02e4", x"02e4", x"02e4", x"02e4", x"02e4", x"02e4", x"02e5", x"02e5", x"02e5", x"02e5", x"02e5", x"02e5", x"02e5", x"02e6", x"02e6", x"02e6", x"02e6", x"02e6", x"02e6", x"02e7", x"02e7", x"02e7", x"02e7", x"02e7", x"02e7", x"02e7", x"02e8", x"02e8", x"02e8", x"02e8", x"02e8", x"02e8", x"02e8", x"02e9", x"02e9", x"02e9", x"02e9", x"02e9", x"02e9", x"02e9", x"02ea", x"02ea", x"02ea", x"02ea", x"02ea", x"02ea", x"02eb", x"02eb", x"02eb", x"02eb", x"02eb", x"02eb", x"02eb", x"02ec", x"02ec", x"02ec", x"02ec", x"02ec", x"02ec", x"02ec", x"02ed", x"02ed", x"02ed", x"02ed", x"02ed", x"02ed", x"02ee", x"02ee", x"02ee", x"02ee", x"02ee", x"02ee", x"02ee", x"02ef", x"02ef", x"02ef", x"02ef", x"02ef", x"02ef", x"02ef", x"02f0", x"02f0", x"02f0", x"02f0", x"02f0", x"02f0", x"02f1", x"02f1", x"02f1", x"02f1", x"02f1", x"02f1", x"02f1", x"02f2", x"02f2", x"02f2", x"02f2", x"02f2", x"02f2", x"02f2", x"02f3", x"02f3", x"02f3", x"02f3", x"02f3", x"02f3", x"02f4", x"02f4", x"02f4", x"02f4", x"02f4", x"02f4", x"02f4", x"02f5", x"02f5", x"02f5", x"02f5", x"02f5", x"02f5", x"02f5", x"02f6", x"02f6", x"02f6", x"02f6", x"02f6", x"02f6", x"02f7", x"02f7", x"02f7", x"02f7", x"02f7", x"02f7", x"02f7", x"02f8", x"02f8", x"02f8", x"02f8", x"02f8", x"02f8", x"02f8", x"02f9", x"02f9", x"02f9", x"02f9", x"02f9", x"02f9", x"02fa", x"02fa", x"02fa", x"02fa", x"02fa", x"02fa", x"02fa", x"02fb", x"02fb", x"02fb", x"02fb", x"02fb", x"02fb", x"02fc", x"02fc", x"02fc", x"02fc", x"02fc", x"02fc", x"02fc", x"02fd", x"02fd", x"02fd", x"02fd", x"02fd", x"02fd", x"02fe", x"02fe", x"02fe", x"02fe", x"02fe", x"02fe", x"02fe", x"02ff", x"02ff", x"02ff", x"02ff", x"02ff", x"02ff", x"02ff", x"0300", x"0300", x"0300", x"0300", x"0300", x"0300", x"0301", x"0301", x"0301", x"0301", x"0301", x"0301", x"0301", x"0302", x"0302", x"0302", x"0302", x"0302", x"0302", x"0303", x"0303", x"0303", x"0303", x"0303", x"0303", x"0303", x"0304", x"0304", x"0304", x"0304", x"0304", x"0304", x"0305", x"0305", x"0305", x"0305", x"0305", x"0305", x"0305", x"0306", x"0306", x"0306", x"0306", x"0306", x"0306", x"0307", x"0307", x"0307", x"0307", x"0307", x"0307", x"0307", x"0308", x"0308", x"0308", x"0308", x"0308", x"0308", x"0309", x"0309", x"0309", x"0309", x"0309", x"0309", x"0309", x"030a", x"030a", x"030a", x"030a", x"030a", x"030a", x"030b", x"030b", x"030b", x"030b", x"030b", x"030b", x"030b", x"030c", x"030c", x"030c", x"030c", x"030c", x"030c", x"030d", x"030d", x"030d", x"030d", x"030d", x"030d", x"030d", x"030e", x"030e", x"030e", x"030e", x"030e", x"030e", x"030f", x"030f", x"030f", x"030f", x"030f", x"030f", x"030f", x"0310", x"0310", x"0310", x"0310", x"0310", x"0310", x"0311", x"0311", x"0311", x"0311", x"0311", x"0311", x"0311", x"0312", x"0312", x"0312", x"0312", x"0312", x"0312", x"0313", x"0313", x"0313", x"0313", x"0313", x"0313", x"0313", x"0314", x"0314", x"0314", x"0314", x"0314", x"0314", x"0315", x"0315", x"0315", x"0315", x"0315", x"0315", x"0316", x"0316", x"0316", x"0316", x"0316", x"0316", x"0316", x"0317", x"0317", x"0317", x"0317", x"0317", x"0317", x"0318", x"0318", x"0318", x"0318", x"0318", x"0318", x"0318", x"0319", x"0319", x"0319", x"0319", x"0319", x"0319", x"031a", x"031a", x"031a", x"031a", x"031a", x"031a", x"031a", x"031b", x"031b", x"031b", x"031b", x"031b", x"031b", x"031c", x"031c", x"031c", x"031c", x"031c", x"031c", x"031d", x"031d", x"031d", x"031d", x"031d", x"031d", x"031d", x"031e", x"031e", x"031e", x"031e", x"031e", x"031e", x"031f", x"031f", x"031f", x"031f", x"031f", x"031f", x"0320", x"0320", x"0320", x"0320", x"0320", x"0320", x"0320", x"0321", x"0321", x"0321", x"0321", x"0321", x"0321", x"0322", x"0322", x"0322", x"0322", x"0322", x"0322", x"0323", x"0323", x"0323", x"0323", x"0323", x"0323", x"0323", x"0324", x"0324", x"0324", x"0324", x"0324", x"0324", x"0325", x"0325", x"0325", x"0325", x"0325", x"0325", x"0326", x"0326", x"0326", x"0326", x"0326", x"0326", x"0326", x"0327", x"0327", x"0327", x"0327", x"0327", x"0327", x"0328", x"0328", x"0328", x"0328", x"0328", x"0328", x"0329", x"0329", x"0329", x"0329", x"0329", x"0329", x"0329", x"032a", x"032a", x"032a", x"032a", x"032a", x"032a", x"032b", x"032b", x"032b", x"032b", x"032b", x"032b", x"032c", x"032c", x"032c", x"032c", x"032c", x"032c", x"032c", x"032d", x"032d", x"032d", x"032d", x"032d", x"032d", x"032e", x"032e", x"032e", x"032e", x"032e", x"032e", x"032f", x"032f", x"032f", x"032f", x"032f", x"032f", x"0330", x"0330", x"0330", x"0330", x"0330", x"0330", x"0330", x"0331", x"0331", x"0331", x"0331", x"0331", x"0331", x"0332", x"0332", x"0332", x"0332", x"0332", x"0332", x"0333", x"0333", x"0333", x"0333", x"0333", x"0333", x"0334", x"0334", x"0334", x"0334", x"0334", x"0334", x"0334", x"0335", x"0335", x"0335", x"0335", x"0335", x"0335", x"0336", x"0336", x"0336", x"0336", x"0336", x"0336", x"0337", x"0337", x"0337", x"0337", x"0337", x"0337", x"0338", x"0338", x"0338", x"0338", x"0338", x"0338", x"0338", x"0339", x"0339", x"0339", x"0339", x"0339", x"0339", x"033a", x"033a", x"033a", x"033a", x"033a", x"033a", x"033b", x"033b", x"033b", x"033b", x"033b", x"033b", x"033c", x"033c", x"033c", x"033c", x"033c", x"033c", x"033d", x"033d", x"033d", x"033d", x"033d", x"033d", x"033d", x"033e", x"033e", x"033e", x"033e", x"033e", x"033e", x"033f", x"033f", x"033f", x"033f", x"033f", x"033f", x"0340", x"0340", x"0340", x"0340", x"0340", x"0340", x"0341", x"0341", x"0341", x"0341", x"0341", x"0341", x"0342", x"0342", x"0342", x"0342", x"0342", x"0342", x"0342", x"0343", x"0343", x"0343", x"0343", x"0343", x"0343", x"0344", x"0344", x"0344", x"0344", x"0344", x"0344", x"0345", x"0345", x"0345", x"0345", x"0345", x"0345", x"0346", x"0346", x"0346", x"0346", x"0346", x"0346", x"0347", x"0347", x"0347", x"0347", x"0347", x"0347", x"0348", x"0348", x"0348", x"0348", x"0348", x"0348", x"0349", x"0349", x"0349", x"0349", x"0349", x"0349", x"0349", x"034a", x"034a", x"034a", x"034a", x"034a", x"034a", x"034b", x"034b", x"034b", x"034b", x"034b", x"034b", x"034c", x"034c", x"034c", x"034c", x"034c", x"034c", x"034d", x"034d", x"034d", x"034d", x"034d", x"034d", x"034e", x"034e", x"034e", x"034e", x"034e", x"034e", x"034f", x"034f", x"034f", x"034f", x"034f", x"034f", x"0350", x"0350", x"0350", x"0350", x"0350", x"0350", x"0351", x"0351", x"0351", x"0351", x"0351", x"0351", x"0352", x"0352", x"0352", x"0352", x"0352", x"0352", x"0353", x"0353", x"0353", x"0353", x"0353", x"0353", x"0353", x"0354", x"0354", x"0354", x"0354", x"0354", x"0354", x"0355", x"0355", x"0355", x"0355", x"0355", x"0355", x"0356", x"0356", x"0356", x"0356", x"0356", x"0356", x"0357", x"0357", x"0357", x"0357", x"0357", x"0357", x"0358", x"0358", x"0358", x"0358", x"0358", x"0358", x"0359", x"0359", x"0359", x"0359", x"0359", x"0359", x"035a", x"035a", x"035a", x"035a", x"035a", x"035a", x"035b", x"035b", x"035b", x"035b", x"035b", x"035b", x"035c", x"035c", x"035c", x"035c", x"035c", x"035c", x"035d", x"035d", x"035d", x"035d", x"035d", x"035d", x"035e", x"035e", x"035e", x"035e", x"035e", x"035e", x"035f", x"035f", x"035f", x"035f", x"035f", x"035f", x"0360", x"0360", x"0360", x"0360", x"0360", x"0360", x"0361", x"0361", x"0361", x"0361", x"0361", x"0361", x"0362", x"0362", x"0362", x"0362", x"0362", x"0362", x"0363", x"0363", x"0363", x"0363", x"0363", x"0363", x"0364", x"0364", x"0364", x"0364", x"0364", x"0364", x"0365", x"0365", x"0365", x"0365", x"0365", x"0365", x"0366", x"0366", x"0366", x"0366", x"0366", x"0366", x"0367", x"0367", x"0367", x"0367", x"0367", x"0367", x"0368", x"0368", x"0368", x"0368", x"0368", x"0368", x"0369", x"0369", x"0369", x"0369", x"0369", x"0369", x"036a", x"036a", x"036a", x"036a", x"036a", x"036a", x"036b", x"036b", x"036b", x"036b", x"036b", x"036b", x"036c", x"036c", x"036c", x"036c", x"036c", x"036c", x"036d", x"036d", x"036d", x"036d", x"036d", x"036d", x"036e", x"036e", x"036e", x"036e", x"036e", x"036e", x"036f", x"036f", x"036f", x"036f", x"036f", x"0370", x"0370", x"0370", x"0370", x"0370", x"0370", x"0371", x"0371", x"0371", x"0371", x"0371", x"0371", x"0372", x"0372", x"0372", x"0372", x"0372", x"0372", x"0373", x"0373", x"0373", x"0373", x"0373", x"0373", x"0374", x"0374", x"0374", x"0374", x"0374", x"0374", x"0375", x"0375", x"0375", x"0375", x"0375", x"0375", x"0376", x"0376", x"0376", x"0376", x"0376", x"0376", x"0377", x"0377", x"0377", x"0377", x"0377", x"0377", x"0378", x"0378", x"0378", x"0378", x"0378", x"0378", x"0379", x"0379", x"0379", x"0379", x"0379", x"0379", x"037a", x"037a", x"037a", x"037a", x"037a", x"037b", x"037b", x"037b", x"037b", x"037b", x"037b", x"037c", x"037c", x"037c", x"037c", x"037c", x"037c", x"037d", x"037d", x"037d", x"037d", x"037d", x"037d", x"037e", x"037e", x"037e", x"037e", x"037e", x"037e", x"037f", x"037f", x"037f", x"037f", x"037f", x"037f", x"0380", x"0380", x"0380", x"0380", x"0380", x"0380", x"0381", x"0381", x"0381", x"0381", x"0381", x"0382", x"0382", x"0382", x"0382", x"0382", x"0382", x"0383", x"0383", x"0383", x"0383", x"0383", x"0383", x"0384", x"0384", x"0384", x"0384", x"0384", x"0384", x"0385", x"0385", x"0385", x"0385", x"0385", x"0385", x"0386", x"0386", x"0386", x"0386", x"0386", x"0386", x"0387", x"0387", x"0387", x"0387", x"0387", x"0388", x"0388", x"0388", x"0388", x"0388", x"0388", x"0389", x"0389", x"0389", x"0389", x"0389", x"0389", x"038a", x"038a", x"038a", x"038a", x"038a", x"038a", x"038b", x"038b", x"038b", x"038b", x"038b", x"038b", x"038c", x"038c", x"038c", x"038c", x"038c", x"038d", x"038d", x"038d", x"038d", x"038d", x"038d", x"038e", x"038e", x"038e", x"038e", x"038e", x"038e", x"038f", x"038f", x"038f", x"038f", x"038f", x"038f", x"0390", x"0390", x"0390", x"0390", x"0390", x"0390", x"0391", x"0391", x"0391", x"0391", x"0391", x"0392", x"0392", x"0392", x"0392", x"0392", x"0392", x"0393", x"0393", x"0393", x"0393", x"0393", x"0393", x"0394", x"0394", x"0394", x"0394", x"0394", x"0394", x"0395", x"0395", x"0395", x"0395", x"0395", x"0396", x"0396", x"0396", x"0396", x"0396", x"0396", x"0397", x"0397", x"0397", x"0397", x"0397", x"0397", x"0398", x"0398", x"0398", x"0398", x"0398", x"0398", x"0399", x"0399", x"0399", x"0399", x"0399", x"039a", x"039a", x"039a", x"039a", x"039a", x"039a", x"039b", x"039b", x"039b", x"039b", x"039b", x"039b", x"039c", x"039c", x"039c", x"039c", x"039c", x"039d", x"039d", x"039d", x"039d", x"039d", x"039d", x"039e", x"039e", x"039e", x"039e", x"039e", x"039e", x"039f", x"039f", x"039f", x"039f", x"039f", x"039f", x"03a0", x"03a0", x"03a0", x"03a0", x"03a0", x"03a1", x"03a1", x"03a1", x"03a1", x"03a1", x"03a1", x"03a2", x"03a2", x"03a2", x"03a2", x"03a2", x"03a2", x"03a3", x"03a3", x"03a3", x"03a3", x"03a3", x"03a4", x"03a4", x"03a4", x"03a4", x"03a4", x"03a4", x"03a5", x"03a5", x"03a5", x"03a5", x"03a5", x"03a5", x"03a6", x"03a6", x"03a6", x"03a6", x"03a6", x"03a7", x"03a7", x"03a7", x"03a7", x"03a7", x"03a7", x"03a8", x"03a8", x"03a8", x"03a8", x"03a8", x"03a8", x"03a9", x"03a9", x"03a9", x"03a9", x"03a9", x"03aa", x"03aa", x"03aa", x"03aa", x"03aa", x"03aa", x"03ab", x"03ab", x"03ab", x"03ab", x"03ab", x"03ab", x"03ac", x"03ac", x"03ac", x"03ac", x"03ac", x"03ad", x"03ad", x"03ad", x"03ad", x"03ad", x"03ad", x"03ae", x"03ae", x"03ae", x"03ae", x"03ae", x"03ae", x"03af", x"03af", x"03af", x"03af", x"03af", x"03b0", x"03b0", x"03b0", x"03b0", x"03b0", x"03b0", x"03b1", x"03b1", x"03b1", x"03b1", x"03b1", x"03b1", x"03b2", x"03b2", x"03b2", x"03b2", x"03b2", x"03b3", x"03b3", x"03b3", x"03b3", x"03b3", x"03b3", x"03b4", x"03b4", x"03b4", x"03b4", x"03b4", x"03b4", x"03b5", x"03b5", x"03b5", x"03b5", x"03b5", x"03b6", x"03b6", x"03b6", x"03b6", x"03b6", x"03b6", x"03b7", x"03b7", x"03b7", x"03b7", x"03b7", x"03b8", x"03b8", x"03b8", x"03b8", x"03b8", x"03b8", x"03b9", x"03b9", x"03b9", x"03b9", x"03b9", x"03b9", x"03ba", x"03ba", x"03ba", x"03ba", x"03ba", x"03bb", x"03bb", x"03bb", x"03bb", x"03bb", x"03bb", x"03bc", x"03bc", x"03bc", x"03bc", x"03bc", x"03bd", x"03bd", x"03bd", x"03bd", x"03bd", x"03bd", x"03be", x"03be", x"03be", x"03be", x"03be", x"03be", x"03bf", x"03bf", x"03bf", x"03bf", x"03bf", x"03c0", x"03c0", x"03c0", x"03c0", x"03c0", x"03c0", x"03c1", x"03c1", x"03c1", x"03c1", x"03c1", x"03c2", x"03c2", x"03c2", x"03c2", x"03c2", x"03c2", x"03c3", x"03c3", x"03c3", x"03c3", x"03c3", x"03c4", x"03c4", x"03c4", x"03c4", x"03c4", x"03c4", x"03c5", x"03c5", x"03c5", x"03c5", x"03c5", x"03c6", x"03c6", x"03c6", x"03c6", x"03c6", x"03c6", x"03c7", x"03c7", x"03c7", x"03c7", x"03c7", x"03c7", x"03c8", x"03c8", x"03c8", x"03c8", x"03c8", x"03c9", x"03c9", x"03c9", x"03c9", x"03c9", x"03c9", x"03ca", x"03ca", x"03ca", x"03ca", x"03ca", x"03cb", x"03cb", x"03cb", x"03cb", x"03cb", x"03cb", x"03cc", x"03cc", x"03cc", x"03cc", x"03cc", x"03cd", x"03cd", x"03cd", x"03cd", x"03cd", x"03cd", x"03ce", x"03ce", x"03ce", x"03ce", x"03ce", x"03cf", x"03cf", x"03cf", x"03cf", x"03cf", x"03cf", x"03d0", x"03d0", x"03d0", x"03d0", x"03d0", x"03d1", x"03d1", x"03d1", x"03d1", x"03d1", x"03d1", x"03d2", x"03d2", x"03d2", x"03d2", x"03d2", x"03d3", x"03d3", x"03d3", x"03d3", x"03d3", x"03d3", x"03d4", x"03d4", x"03d4", x"03d4", x"03d4", x"03d5", x"03d5", x"03d5", x"03d5", x"03d5", x"03d5", x"03d6", x"03d6", x"03d6", x"03d6", x"03d6", x"03d7", x"03d7", x"03d7", x"03d7", x"03d7", x"03d7", x"03d8", x"03d8", x"03d8", x"03d8", x"03d8", x"03d9", x"03d9", x"03d9", x"03d9", x"03d9", x"03d9", x"03da", x"03da", x"03da", x"03da", x"03da", x"03db", x"03db", x"03db", x"03db", x"03db", x"03db", x"03dc", x"03dc", x"03dc", x"03dc", x"03dc", x"03dd", x"03dd", x"03dd", x"03dd", x"03dd", x"03dd", x"03de", x"03de", x"03de", x"03de", x"03de", x"03df", x"03df", x"03df", x"03df", x"03df", x"03e0", x"03e0", x"03e0", x"03e0", x"03e0", x"03e0", x"03e1", x"03e1", x"03e1", x"03e1", x"03e1", x"03e2", x"03e2", x"03e2", x"03e2", x"03e2", x"03e2", x"03e3", x"03e3", x"03e3", x"03e3", x"03e3", x"03e4", x"03e4", x"03e4", x"03e4", x"03e4", x"03e4", x"03e5", x"03e5", x"03e5", x"03e5", x"03e5", x"03e6", x"03e6", x"03e6", x"03e6", x"03e6", x"03e7", x"03e7", x"03e7", x"03e7", x"03e7", x"03e7", x"03e8", x"03e8", x"03e8", x"03e8", x"03e8", x"03e9", x"03e9", x"03e9", x"03e9", x"03e9", x"03e9", x"03ea", x"03ea", x"03ea", x"03ea", x"03ea", x"03eb", x"03eb", x"03eb", x"03eb", x"03eb", x"03eb", x"03ec", x"03ec", x"03ec", x"03ec", x"03ec", x"03ed", x"03ed", x"03ed", x"03ed", x"03ed", x"03ee", x"03ee", x"03ee", x"03ee", x"03ee", x"03ee", x"03ef", x"03ef", x"03ef", x"03ef", x"03ef", x"03f0", x"03f0", x"03f0", x"03f0", x"03f0", x"03f0", x"03f1", x"03f1", x"03f1", x"03f1", x"03f1", x"03f2", x"03f2", x"03f2", x"03f2", x"03f2", x"03f3", x"03f3", x"03f3", x"03f3", x"03f3", x"03f3", x"03f4", x"03f4", x"03f4", x"03f4", x"03f4", x"03f5", x"03f5", x"03f5", x"03f5", x"03f5", x"03f6", x"03f6", x"03f6", x"03f6", x"03f6", x"03f6", x"03f7", x"03f7", x"03f7", x"03f7", x"03f7", x"03f8", x"03f8", x"03f8", x"03f8", x"03f8", x"03f9", x"03f9", x"03f9", x"03f9", x"03f9", x"03f9", x"03fa", x"03fa", x"03fa", x"03fa", x"03fa", x"03fb", x"03fb", x"03fb", x"03fb", x"03fb", x"03fb", x"03fc", x"03fc", x"03fc", x"03fc", x"03fc", x"03fd", x"03fd", x"03fd", x"03fd", x"03fd", x"03fe", x"03fe", x"03fe", x"03fe", x"03fe", x"03fe", x"03ff", x"03ff", x"03ff", x"03ff", x"03ff", x"0400", x"0400", x"0400", x"0400", x"0400", x"0401", x"0401", x"0401", x"0401", x"0401", x"0401", x"0402", x"0402", x"0402", x"0402", x"0402", x"0403", x"0403", x"0403", x"0403", x"0403", x"0404", x"0404", x"0404", x"0404", x"0404", x"0404", x"0405", x"0405", x"0405", x"0405", x"0405", x"0406", x"0406", x"0406", x"0406", x"0406", x"0407", x"0407", x"0407", x"0407", x"0407", x"0408", x"0408", x"0408", x"0408", x"0408", x"0408", x"0409", x"0409", x"0409", x"0409", x"0409", x"040a", x"040a", x"040a", x"040a", x"040a", x"040b", x"040b", x"040b", x"040b", x"040b", x"040b", x"040c", x"040c", x"040c", x"040c", x"040c", x"040d", x"040d", x"040d", x"040d", x"040d", x"040e", x"040e", x"040e", x"040e", x"040e", x"040e", x"040f", x"040f", x"040f", x"040f", x"040f", x"0410", x"0410", x"0410", x"0410", x"0410", x"0411", x"0411", x"0411", x"0411", x"0411", x"0412", x"0412", x"0412", x"0412", x"0412", x"0412", x"0413", x"0413", x"0413", x"0413", x"0413", x"0414", x"0414", x"0414", x"0414", x"0414", x"0415", x"0415", x"0415", x"0415", x"0415", x"0416", x"0416", x"0416", x"0416", x"0416", x"0416", x"0417", x"0417", x"0417", x"0417", x"0417", x"0418", x"0418", x"0418", x"0418", x"0418", x"0419", x"0419", x"0419", x"0419", x"0419", x"041a", x"041a", x"041a", x"041a", x"041a", x"041a", x"041b", x"041b", x"041b", x"041b", x"041b", x"041c", x"041c", x"041c", x"041c", x"041c", x"041d", x"041d", x"041d", x"041d", x"041d", x"041e", x"041e", x"041e", x"041e", x"041e", x"041e", x"041f", x"041f", x"041f", x"041f", x"041f", x"0420", x"0420", x"0420", x"0420", x"0420", x"0421", x"0421", x"0421", x"0421", x"0421", x"0422", x"0422", x"0422", x"0422", x"0422", x"0422", x"0423", x"0423", x"0423", x"0423", x"0423", x"0424", x"0424", x"0424", x"0424", x"0424", x"0425", x"0425", x"0425", x"0425", x"0425", x"0426", x"0426", x"0426", x"0426", x"0426", x"0427", x"0427", x"0427", x"0427", x"0427", x"0427", x"0428", x"0428", x"0428", x"0428", x"0428", x"0429", x"0429", x"0429", x"0429", x"0429", x"042a", x"042a", x"042a", x"042a", x"042a", x"042b", x"042b", x"042b", x"042b", x"042b", x"042c", x"042c", x"042c", x"042c", x"042c", x"042c", x"042d", x"042d", x"042d", x"042d", x"042d", x"042e", x"042e", x"042e", x"042e", x"042e", x"042f", x"042f", x"042f", x"042f", x"042f", x"0430", x"0430", x"0430", x"0430", x"0430", x"0431", x"0431", x"0431", x"0431", x"0431", x"0432", x"0432", x"0432", x"0432", x"0432", x"0432", x"0433", x"0433", x"0433", x"0433", x"0433", x"0434", x"0434", x"0434", x"0434", x"0434", x"0435", x"0435", x"0435", x"0435", x"0435", x"0436", x"0436", x"0436", x"0436", x"0436", x"0437", x"0437", x"0437", x"0437", x"0437", x"0438", x"0438", x"0438", x"0438", x"0438", x"0438", x"0439", x"0439", x"0439", x"0439", x"0439", x"043a", x"043a", x"043a", x"043a", x"043a", x"043b", x"043b", x"043b", x"043b", x"043b", x"043c", x"043c", x"043c", x"043c", x"043c", x"043d", x"043d", x"043d", x"043d", x"043d", x"043e", x"043e", x"043e", x"043e", x"043e", x"043f", x"043f", x"043f", x"043f", x"043f", x"0440", x"0440", x"0440", x"0440", x"0440", x"0440", x"0441", x"0441", x"0441", x"0441", x"0441", x"0442", x"0442", x"0442", x"0442", x"0442", x"0443", x"0443", x"0443", x"0443", x"0443", x"0444", x"0444", x"0444", x"0444", x"0444", x"0445", x"0445", x"0445", x"0445", x"0445", x"0446", x"0446", x"0446", x"0446", x"0446", x"0447", x"0447", x"0447", x"0447", x"0447", x"0448", x"0448", x"0448", x"0448", x"0448", x"0448", x"0449", x"0449", x"0449", x"0449", x"0449", x"044a", x"044a", x"044a", x"044a", x"044a", x"044b", x"044b", x"044b", x"044b", x"044b", x"044c", x"044c", x"044c", x"044c", x"044c", x"044d", x"044d", x"044d", x"044d", x"044d", x"044e", x"044e", x"044e", x"044e", x"044e", x"044f", x"044f", x"044f", x"044f", x"044f", x"0450", x"0450", x"0450", x"0450", x"0450", x"0451", x"0451", x"0451", x"0451", x"0451", x"0452", x"0452", x"0452", x"0452", x"0452", x"0453", x"0453", x"0453", x"0453", x"0453", x"0454", x"0454", x"0454", x"0454", x"0454", x"0454", x"0455", x"0455", x"0455", x"0455", x"0455", x"0456", x"0456", x"0456", x"0456", x"0456", x"0457", x"0457", x"0457", x"0457", x"0457", x"0458", x"0458", x"0458", x"0458", x"0458", x"0459", x"0459", x"0459", x"0459", x"0459", x"045a", x"045a", x"045a", x"045a", x"045a", x"045b", x"045b", x"045b", x"045b", x"045b", x"045c", x"045c", x"045c", x"045c", x"045c", x"045d", x"045d", x"045d", x"045d", x"045d", x"045e", x"045e", x"045e", x"045e", x"045e", x"045f", x"045f", x"045f", x"045f", x"045f", x"0460", x"0460", x"0460", x"0460", x"0460", x"0461", x"0461", x"0461", x"0461", x"0461", x"0462", x"0462", x"0462", x"0462", x"0462", x"0463", x"0463", x"0463", x"0463", x"0463", x"0464", x"0464", x"0464", x"0464", x"0464", x"0465", x"0465", x"0465", x"0465", x"0465", x"0466", x"0466", x"0466", x"0466", x"0466", x"0467", x"0467", x"0467", x"0467", x"0467", x"0468", x"0468", x"0468", x"0468", x"0468", x"0469", x"0469", x"0469", x"0469", x"0469", x"046a", x"046a", x"046a", x"046a", x"046a", x"046b", x"046b", x"046b", x"046b", x"046b", x"046c", x"046c", x"046c", x"046c", x"046c", x"046d", x"046d", x"046d", x"046d", x"046d", x"046e", x"046e", x"046e", x"046e", x"046e", x"046f", x"046f", x"046f", x"046f", x"046f", x"0470", x"0470", x"0470", x"0470", x"0470", x"0471", x"0471", x"0471", x"0471", x"0471", x"0472", x"0472", x"0472", x"0472", x"0472", x"0473", x"0473", x"0473", x"0473", x"0473", x"0474", x"0474", x"0474", x"0474", x"0474", x"0475", x"0475", x"0475", x"0475", x"0475", x"0476", x"0476", x"0476", x"0476", x"0476", x"0477", x"0477", x"0477", x"0477", x"0477", x"0478", x"0478", x"0478", x"0478", x"0478", x"0479", x"0479", x"0479", x"0479", x"0479", x"047a", x"047a", x"047a", x"047a", x"047a", x"047b", x"047b", x"047b", x"047b", x"047b", x"047c", x"047c", x"047c", x"047c", x"047c", x"047d", x"047d", x"047d", x"047d", x"047d", x"047e", x"047e", x"047e", x"047e", x"047e", x"047f", x"047f", x"047f", x"047f", x"047f", x"0480", x"0480", x"0480", x"0480", x"0480", x"0481", x"0481", x"0481", x"0481", x"0481", x"0482", x"0482", x"0482", x"0482", x"0482", x"0483", x"0483", x"0483", x"0483", x"0483", x"0484", x"0484", x"0484", x"0484", x"0485", x"0485", x"0485", x"0485", x"0485", x"0486", x"0486", x"0486", x"0486", x"0486", x"0487", x"0487", x"0487", x"0487", x"0487", x"0488", x"0488", x"0488", x"0488", x"0488", x"0489", x"0489", x"0489", x"0489", x"0489", x"048a", x"048a", x"048a", x"048a", x"048a", x"048b", x"048b", x"048b", x"048b", x"048b", x"048c", x"048c", x"048c", x"048c", x"048c", x"048d", x"048d", x"048d", x"048d", x"048d", x"048e", x"048e", x"048e", x"048e", x"048e", x"048f", x"048f", x"048f", x"048f", x"048f", x"0490", x"0490", x"0490", x"0490", x"0491", x"0491", x"0491", x"0491", x"0491", x"0492", x"0492", x"0492", x"0492", x"0492", x"0493", x"0493", x"0493", x"0493", x"0493", x"0494", x"0494", x"0494", x"0494", x"0494", x"0495", x"0495", x"0495", x"0495", x"0495", x"0496", x"0496", x"0496", x"0496", x"0496", x"0497", x"0497", x"0497", x"0497", x"0497", x"0498", x"0498", x"0498", x"0498", x"0498", x"0499", x"0499", x"0499", x"0499", x"0499", x"049a", x"049a", x"049a", x"049a", x"049b", x"049b", x"049b", x"049b", x"049b", x"049c", x"049c", x"049c", x"049c", x"049c", x"049d", x"049d", x"049d", x"049d", x"049d", x"049e", x"049e", x"049e", x"049e", x"049e", x"049f", x"049f", x"049f", x"049f", x"049f", x"04a0", x"04a0", x"04a0", x"04a0", x"04a0", x"04a1", x"04a1", x"04a1", x"04a1", x"04a2", x"04a2", x"04a2", x"04a2", x"04a2", x"04a3", x"04a3", x"04a3", x"04a3", x"04a3", x"04a4", x"04a4", x"04a4", x"04a4", x"04a4", x"04a5", x"04a5", x"04a5", x"04a5", x"04a5", x"04a6", x"04a6", x"04a6", x"04a6", x"04a6", x"04a7", x"04a7", x"04a7", x"04a7", x"04a7", x"04a8", x"04a8", x"04a8", x"04a8", x"04a9", x"04a9", x"04a9", x"04a9", x"04a9", x"04aa", x"04aa", x"04aa", x"04aa", x"04aa", x"04ab", x"04ab", x"04ab", x"04ab", x"04ab", x"04ac", x"04ac", x"04ac", x"04ac", x"04ac", x"04ad", x"04ad", x"04ad", x"04ad", x"04ad", x"04ae", x"04ae", x"04ae", x"04ae", x"04af", x"04af", x"04af", x"04af", x"04af", x"04b0", x"04b0", x"04b0", x"04b0", x"04b0", x"04b1", x"04b1", x"04b1", x"04b1", x"04b1", x"04b2", x"04b2", x"04b2", x"04b2", x"04b2", x"04b3", x"04b3", x"04b3", x"04b3", x"04b3", x"04b4", x"04b4", x"04b4", x"04b4", x"04b5", x"04b5", x"04b5", x"04b5", x"04b5", x"04b6", x"04b6", x"04b6", x"04b6", x"04b6", x"04b7", x"04b7", x"04b7", x"04b7", x"04b7", x"04b8", x"04b8", x"04b8", x"04b8", x"04b8", x"04b9", x"04b9", x"04b9", x"04b9", x"04ba", x"04ba", x"04ba", x"04ba", x"04ba", x"04bb", x"04bb", x"04bb", x"04bb", x"04bb", x"04bc", x"04bc", x"04bc", x"04bc", x"04bc", x"04bd", x"04bd", x"04bd", x"04bd", x"04bd", x"04be", x"04be", x"04be", x"04be", x"04bf", x"04bf", x"04bf", x"04bf", x"04bf", x"04c0", x"04c0", x"04c0", x"04c0", x"04c0", x"04c1", x"04c1", x"04c1", x"04c1", x"04c1", x"04c2", x"04c2", x"04c2", x"04c2", x"04c2", x"04c3", x"04c3", x"04c3", x"04c3", x"04c4", x"04c4", x"04c4", x"04c4", x"04c4", x"04c5", x"04c5", x"04c5", x"04c5", x"04c5", x"04c6", x"04c6", x"04c6", x"04c6", x"04c6", x"04c7", x"04c7", x"04c7", x"04c7", x"04c7", x"04c8", x"04c8", x"04c8", x"04c8", x"04c9", x"04c9", x"04c9", x"04c9", x"04c9", x"04ca", x"04ca", x"04ca", x"04ca", x"04ca", x"04cb", x"04cb", x"04cb", x"04cb", x"04cb", x"04cc", x"04cc", x"04cc", x"04cc", x"04cd", x"04cd", x"04cd", x"04cd", x"04cd", x"04ce", x"04ce", x"04ce", x"04ce", x"04ce", x"04cf", x"04cf", x"04cf", x"04cf", x"04cf", x"04d0", x"04d0", x"04d0", x"04d0", x"04d1", x"04d1", x"04d1", x"04d1", x"04d1", x"04d2", x"04d2", x"04d2", x"04d2", x"04d2", x"04d3", x"04d3", x"04d3", x"04d3", x"04d3", x"04d4", x"04d4", x"04d4", x"04d4", x"04d5", x"04d5", x"04d5", x"04d5", x"04d5", x"04d6", x"04d6", x"04d6", x"04d6", x"04d6", x"04d7", x"04d7", x"04d7", x"04d7", x"04d7", x"04d8", x"04d8", x"04d8", x"04d8", x"04d9", x"04d9", x"04d9", x"04d9", x"04d9", x"04da", x"04da", x"04da", x"04da", x"04da", x"04db", x"04db", x"04db", x"04db", x"04db", x"04dc", x"04dc", x"04dc", x"04dc", x"04dd", x"04dd", x"04dd", x"04dd", x"04dd", x"04de", x"04de", x"04de", x"04de", x"04de", x"04df", x"04df", x"04df", x"04df", x"04e0", x"04e0", x"04e0", x"04e0", x"04e0", x"04e1", x"04e1", x"04e1", x"04e1", x"04e1", x"04e2", x"04e2", x"04e2", x"04e2", x"04e2", x"04e3", x"04e3", x"04e3", x"04e3", x"04e4", x"04e4", x"04e4", x"04e4", x"04e4", x"04e5", x"04e5", x"04e5", x"04e5", x"04e5", x"04e6", x"04e6", x"04e6", x"04e6", x"04e7", x"04e7", x"04e7", x"04e7", x"04e7", x"04e8", x"04e8", x"04e8", x"04e8", x"04e8", x"04e9", x"04e9", x"04e9", x"04e9", x"04e9", x"04ea", x"04ea", x"04ea", x"04ea", x"04eb", x"04eb", x"04eb", x"04eb", x"04eb", x"04ec", x"04ec", x"04ec", x"04ec", x"04ec", x"04ed", x"04ed", x"04ed", x"04ed", x"04ee", x"04ee", x"04ee", x"04ee", x"04ee", x"04ef", x"04ef", x"04ef", x"04ef", x"04ef", x"04f0", x"04f0", x"04f0", x"04f0", x"04f1", x"04f1", x"04f1", x"04f1", x"04f1", x"04f2", x"04f2", x"04f2", x"04f2", x"04f2", x"04f3", x"04f3", x"04f3", x"04f3", x"04f4", x"04f4", x"04f4", x"04f4", x"04f4", x"04f5", x"04f5", x"04f5", x"04f5", x"04f5", x"04f6", x"04f6", x"04f6", x"04f6", x"04f7", x"04f7", x"04f7", x"04f7", x"04f7", x"04f8", x"04f8", x"04f8", x"04f8", x"04f8", x"04f9", x"04f9", x"04f9", x"04f9", x"04fa", x"04fa", x"04fa", x"04fa", x"04fa", x"04fb", x"04fb", x"04fb", x"04fb", x"04fb", x"04fc", x"04fc", x"04fc", x"04fc", x"04fd", x"04fd", x"04fd", x"04fd", x"04fd", x"04fe", x"04fe", x"04fe", x"04fe", x"04fe", x"04ff", x"04ff", x"04ff", x"04ff", x"0500", x"0500", x"0500", x"0500", x"0500", x"0501", x"0501", x"0501", x"0501", x"0501", x"0502", x"0502", x"0502", x"0502", x"0503", x"0503", x"0503", x"0503", x"0503", x"0504", x"0504", x"0504", x"0504", x"0504", x"0505", x"0505", x"0505", x"0505", x"0506", x"0506", x"0506", x"0506", x"0506", x"0507", x"0507", x"0507", x"0507", x"0507", x"0508", x"0508", x"0508", x"0508", x"0509", x"0509", x"0509", x"0509", x"0509", x"050a", x"050a", x"050a", x"050a", x"050a", x"050b", x"050b", x"050b", x"050b", x"050c", x"050c", x"050c", x"050c", x"050c", x"050d", x"050d", x"050d", x"050d", x"050e", x"050e", x"050e", x"050e", x"050e", x"050f", x"050f", x"050f", x"050f", x"050f", x"0510", x"0510", x"0510", x"0510", x"0511", x"0511", x"0511", x"0511", x"0511", x"0512", x"0512", x"0512", x"0512", x"0512", x"0513", x"0513", x"0513", x"0513", x"0514", x"0514", x"0514", x"0514", x"0514", x"0515", x"0515", x"0515", x"0515", x"0516", x"0516", x"0516", x"0516", x"0516", x"0517", x"0517", x"0517", x"0517", x"0517", x"0518", x"0518", x"0518", x"0518", x"0519", x"0519", x"0519", x"0519", x"0519", x"051a", x"051a", x"051a", x"051a", x"051b", x"051b", x"051b", x"051b", x"051b", x"051c", x"051c", x"051c", x"051c", x"051c", x"051d", x"051d", x"051d", x"051d", x"051e", x"051e", x"051e", x"051e", x"051e", x"051f", x"051f", x"051f", x"051f", x"0520", x"0520", x"0520", x"0520", x"0520", x"0521", x"0521", x"0521", x"0521", x"0521", x"0522", x"0522", x"0522", x"0522", x"0523", x"0523", x"0523", x"0523", x"0523", x"0524", x"0524", x"0524", x"0524", x"0525", x"0525", x"0525", x"0525", x"0525", x"0526", x"0526", x"0526", x"0526", x"0526", x"0527", x"0527", x"0527", x"0527", x"0528", x"0528", x"0528", x"0528", x"0528", x"0529", x"0529", x"0529", x"0529", x"052a", x"052a", x"052a", x"052a", x"052a", x"052b", x"052b", x"052b", x"052b", x"052c", x"052c", x"052c", x"052c", x"052c", x"052d", x"052d", x"052d", x"052d", x"052d", x"052e", x"052e", x"052e", x"052e", x"052f", x"052f", x"052f", x"052f", x"052f", x"0530", x"0530", x"0530", x"0530", x"0531", x"0531", x"0531", x"0531", x"0531", x"0532", x"0532", x"0532", x"0532", x"0533", x"0533", x"0533", x"0533", x"0533", x"0534", x"0534", x"0534", x"0534", x"0535", x"0535", x"0535", x"0535", x"0535", x"0536", x"0536", x"0536", x"0536", x"0536", x"0537", x"0537", x"0537", x"0537", x"0538", x"0538", x"0538", x"0538", x"0538", x"0539", x"0539", x"0539", x"0539", x"053a", x"053a", x"053a", x"053a", x"053a", x"053b", x"053b", x"053b", x"053b", x"053c", x"053c", x"053c", x"053c", x"053c", x"053d", x"053d", x"053d", x"053d", x"053e", x"053e", x"053e", x"053e", x"053e", x"053f", x"053f", x"053f", x"053f", x"0540", x"0540", x"0540", x"0540", x"0540", x"0541", x"0541", x"0541", x"0541", x"0541", x"0542", x"0542", x"0542", x"0542", x"0543", x"0543", x"0543", x"0543", x"0543", x"0544", x"0544", x"0544", x"0544", x"0545", x"0545", x"0545", x"0545", x"0545", x"0546", x"0546", x"0546", x"0546", x"0547", x"0547", x"0547", x"0547", x"0547", x"0548", x"0548", x"0548", x"0548", x"0549", x"0549", x"0549", x"0549", x"0549", x"054a", x"054a", x"054a", x"054a", x"054b", x"054b", x"054b", x"054b", x"054b", x"054c", x"054c", x"054c", x"054c", x"054d", x"054d", x"054d", x"054d", x"054d", x"054e", x"054e", x"054e", x"054e", x"054f", x"054f", x"054f", x"054f", x"054f", x"0550", x"0550", x"0550", x"0550", x"0551", x"0551", x"0551", x"0551", x"0551", x"0552", x"0552", x"0552", x"0552", x"0553", x"0553", x"0553", x"0553", x"0553", x"0554", x"0554", x"0554", x"0554", x"0555", x"0555", x"0555", x"0555", x"0555", x"0556", x"0556", x"0556", x"0556", x"0557", x"0557", x"0557", x"0557", x"0557", x"0558", x"0558", x"0558", x"0558", x"0559", x"0559", x"0559", x"0559", x"0559", x"055a", x"055a", x"055a", x"055a", x"055b", x"055b", x"055b", x"055b", x"055b", x"055c", x"055c", x"055c", x"055c", x"055d", x"055d", x"055d", x"055d", x"055d", x"055e", x"055e", x"055e", x"055e", x"055f", x"055f", x"055f", x"055f", x"055f", x"0560", x"0560", x"0560", x"0560", x"0561", x"0561", x"0561", x"0561", x"0561", x"0562", x"0562", x"0562", x"0562", x"0563", x"0563", x"0563", x"0563", x"0563", x"0564", x"0564", x"0564", x"0564", x"0565", x"0565", x"0565", x"0565", x"0565", x"0566", x"0566", x"0566", x"0566", x"0567", x"0567", x"0567", x"0567", x"0567", x"0568", x"0568", x"0568", x"0568", x"0569", x"0569", x"0569", x"0569", x"0569", x"056a", x"056a", x"056a", x"056a", x"056b", x"056b", x"056b", x"056b", x"056c", x"056c", x"056c", x"056c", x"056c", x"056d", x"056d", x"056d", x"056d", x"056e", x"056e", x"056e", x"056e", x"056e", x"056f", x"056f", x"056f", x"056f", x"0570", x"0570", x"0570", x"0570", x"0570", x"0571", x"0571", x"0571", x"0571", x"0572", x"0572", x"0572", x"0572", x"0572", x"0573", x"0573", x"0573", x"0573", x"0574", x"0574", x"0574", x"0574", x"0574", x"0575", x"0575", x"0575", x"0575", x"0576", x"0576", x"0576", x"0576", x"0577", x"0577", x"0577", x"0577", x"0577", x"0578", x"0578", x"0578", x"0578", x"0579", x"0579", x"0579", x"0579", x"0579", x"057a", x"057a", x"057a", x"057a", x"057b", x"057b", x"057b", x"057b", x"057b", x"057c", x"057c", x"057c", x"057c", x"057d", x"057d", x"057d", x"057d", x"057d", x"057e", x"057e", x"057e", x"057e", x"057f", x"057f", x"057f", x"057f", x"0580", x"0580", x"0580", x"0580", x"0580", x"0581", x"0581", x"0581", x"0581", x"0582", x"0582", x"0582", x"0582", x"0582", x"0583", x"0583", x"0583", x"0583", x"0584", x"0584", x"0584", x"0584", x"0584", x"0585", x"0585", x"0585", x"0585", x"0586", x"0586", x"0586", x"0586", x"0587", x"0587", x"0587", x"0587", x"0587", x"0588", x"0588", x"0588", x"0588", x"0589", x"0589", x"0589", x"0589", x"0589", x"058a", x"058a", x"058a", x"058a", x"058b", x"058b", x"058b", x"058b", x"058b", x"058c", x"058c", x"058c", x"058c", x"058d", x"058d", x"058d", x"058d", x"058e", x"058e", x"058e", x"058e", x"058e", x"058f", x"058f", x"058f", x"058f", x"0590", x"0590", x"0590", x"0590", x"0590", x"0591", x"0591", x"0591", x"0591", x"0592", x"0592", x"0592", x"0592", x"0593", x"0593", x"0593", x"0593", x"0593", x"0594", x"0594", x"0594", x"0594", x"0595", x"0595", x"0595", x"0595", x"0595", x"0596", x"0596", x"0596", x"0596", x"0597", x"0597", x"0597", x"0597", x"0598", x"0598", x"0598", x"0598", x"0598", x"0599", x"0599", x"0599", x"0599", x"059a", x"059a", x"059a", x"059a", x"059a", x"059b", x"059b", x"059b", x"059b", x"059c", x"059c", x"059c", x"059c", x"059d", x"059d", x"059d", x"059d", x"059d", x"059e", x"059e", x"059e", x"059e", x"059f", x"059f", x"059f", x"059f", x"059f", x"05a0", x"05a0", x"05a0", x"05a0", x"05a1", x"05a1", x"05a1", x"05a1", x"05a2", x"05a2", x"05a2", x"05a2", x"05a2", x"05a3", x"05a3", x"05a3", x"05a3", x"05a4", x"05a4", x"05a4", x"05a4", x"05a5", x"05a5", x"05a5", x"05a5", x"05a5", x"05a6", x"05a6", x"05a6", x"05a6", x"05a7", x"05a7", x"05a7", x"05a7", x"05a7", x"05a8", x"05a8", x"05a8", x"05a8", x"05a9", x"05a9", x"05a9", x"05a9", x"05aa", x"05aa", x"05aa", x"05aa", x"05aa", x"05ab", x"05ab", x"05ab", x"05ab", x"05ac", x"05ac", x"05ac", x"05ac", x"05ad", x"05ad", x"05ad", x"05ad", x"05ad", x"05ae", x"05ae", x"05ae", x"05ae", x"05af", x"05af", x"05af", x"05af", x"05af", x"05b0", x"05b0", x"05b0", x"05b0", x"05b1", x"05b1", x"05b1", x"05b1", x"05b2", x"05b2", x"05b2", x"05b2", x"05b2", x"05b3", x"05b3", x"05b3", x"05b3", x"05b4", x"05b4", x"05b4", x"05b4", x"05b5", x"05b5", x"05b5", x"05b5", x"05b5", x"05b6", x"05b6", x"05b6", x"05b6", x"05b7", x"05b7", x"05b7", x"05b7", x"05b8", x"05b8", x"05b8", x"05b8", x"05b8", x"05b9", x"05b9", x"05b9", x"05b9", x"05ba", x"05ba", x"05ba", x"05ba", x"05ba", x"05bb", x"05bb", x"05bb", x"05bb", x"05bc", x"05bc", x"05bc", x"05bc", x"05bd", x"05bd", x"05bd", x"05bd", x"05bd", x"05be", x"05be", x"05be", x"05be", x"05bf", x"05bf", x"05bf", x"05bf", x"05c0", x"05c0", x"05c0", x"05c0", x"05c0", x"05c1", x"05c1", x"05c1", x"05c1", x"05c2", x"05c2", x"05c2", x"05c2", x"05c3", x"05c3", x"05c3", x"05c3", x"05c3", x"05c4", x"05c4", x"05c4", x"05c4", x"05c5", x"05c5", x"05c5", x"05c5", x"05c6", x"05c6", x"05c6", x"05c6", x"05c6", x"05c7", x"05c7", x"05c7", x"05c7", x"05c8", x"05c8", x"05c8", x"05c8", x"05c9", x"05c9", x"05c9", x"05c9", x"05c9", x"05ca", x"05ca", x"05ca", x"05ca", x"05cb", x"05cb", x"05cb", x"05cb", x"05cc", x"05cc", x"05cc", x"05cc", x"05cc", x"05cd", x"05cd", x"05cd", x"05cd", x"05ce", x"05ce", x"05ce", x"05ce", x"05cf", x"05cf", x"05cf", x"05cf", x"05cf", x"05d0", x"05d0", x"05d0", x"05d0", x"05d1", x"05d1", x"05d1", x"05d1", x"05d2", x"05d2", x"05d2", x"05d2", x"05d2", x"05d3", x"05d3", x"05d3", x"05d3", x"05d4", x"05d4", x"05d4", x"05d4", x"05d5", x"05d5", x"05d5", x"05d5", x"05d5", x"05d6", x"05d6", x"05d6", x"05d6", x"05d7", x"05d7", x"05d7", x"05d7", x"05d8", x"05d8", x"05d8", x"05d8", x"05d9", x"05d9", x"05d9", x"05d9", x"05d9", x"05da", x"05da", x"05da", x"05da", x"05db", x"05db", x"05db", x"05db", x"05dc", x"05dc", x"05dc", x"05dc", x"05dc", x"05dd", x"05dd", x"05dd", x"05dd", x"05de", x"05de", x"05de", x"05de", x"05df", x"05df", x"05df", x"05df", x"05df", x"05e0", x"05e0", x"05e0", x"05e0", x"05e1", x"05e1", x"05e1", x"05e1", x"05e2", x"05e2", x"05e2", x"05e2", x"05e2", x"05e3", x"05e3", x"05e3", x"05e3", x"05e4", x"05e4", x"05e4", x"05e4", x"05e5", x"05e5", x"05e5", x"05e5", x"05e6", x"05e6", x"05e6", x"05e6", x"05e6", x"05e7", x"05e7", x"05e7", x"05e7", x"05e8", x"05e8", x"05e8", x"05e8", x"05e9", x"05e9", x"05e9", x"05e9", x"05e9", x"05ea", x"05ea", x"05ea", x"05ea", x"05eb", x"05eb", x"05eb", x"05eb", x"05ec", x"05ec", x"05ec", x"05ec", x"05ed", x"05ed", x"05ed", x"05ed", x"05ed", x"05ee", x"05ee", x"05ee", x"05ee", x"05ef", x"05ef", x"05ef", x"05ef", x"05f0", x"05f0", x"05f0", x"05f0", x"05f0", x"05f1", x"05f1", x"05f1", x"05f1", x"05f2", x"05f2", x"05f2", x"05f2", x"05f3", x"05f3", x"05f3", x"05f3", x"05f4", x"05f4", x"05f4", x"05f4", x"05f4", x"05f5", x"05f5", x"05f5", x"05f5", x"05f6", x"05f6", x"05f6", x"05f6", x"05f7", x"05f7", x"05f7", x"05f7", x"05f7", x"05f8", x"05f8", x"05f8", x"05f8", x"05f9", x"05f9", x"05f9", x"05f9", x"05fa", x"05fa", x"05fa", x"05fa", x"05fb", x"05fb", x"05fb", x"05fb", x"05fb", x"05fc", x"05fc", x"05fc", x"05fc", x"05fd", x"05fd", x"05fd", x"05fd", x"05fe", x"05fe", x"05fe", x"05fe", x"05ff", x"05ff", x"05ff", x"05ff", x"05ff", x"0600", x"0600", x"0600", x"0600", x"0601", x"0601", x"0601", x"0601", x"0602", x"0602", x"0602", x"0602", x"0602", x"0603", x"0603", x"0603", x"0603", x"0604", x"0604", x"0604", x"0604", x"0605", x"0605", x"0605", x"0605", x"0606", x"0606", x"0606", x"0606", x"0606", x"0607", x"0607", x"0607", x"0607", x"0608", x"0608", x"0608", x"0608", x"0609", x"0609", x"0609", x"0609", x"060a", x"060a", x"060a", x"060a", x"060a", x"060b", x"060b", x"060b", x"060b", x"060c", x"060c", x"060c", x"060c", x"060d", x"060d", x"060d", x"060d", x"060e", x"060e", x"060e", x"060e", x"060e", x"060f", x"060f", x"060f", x"060f", x"0610", x"0610", x"0610", x"0610", x"0611", x"0611", x"0611", x"0611", x"0612", x"0612", x"0612", x"0612", x"0612", x"0613", x"0613", x"0613", x"0613", x"0614", x"0614", x"0614", x"0614", x"0615", x"0615", x"0615", x"0615", x"0616", x"0616", x"0616", x"0616", x"0616", x"0617", x"0617", x"0617", x"0617", x"0618", x"0618", x"0618", x"0618", x"0619", x"0619", x"0619", x"0619", x"061a", x"061a", x"061a", x"061a", x"061a", x"061b", x"061b", x"061b", x"061b", x"061c", x"061c", x"061c", x"061c", x"061d", x"061d", x"061d", x"061d", x"061e", x"061e", x"061e", x"061e", x"061e", x"061f", x"061f", x"061f", x"061f", x"0620", x"0620", x"0620", x"0620", x"0621", x"0621", x"0621", x"0621", x"0622", x"0622", x"0622", x"0622", x"0623", x"0623", x"0623", x"0623", x"0623", x"0624", x"0624", x"0624", x"0624", x"0625", x"0625", x"0625", x"0625", x"0626", x"0626", x"0626", x"0626", x"0627", x"0627", x"0627", x"0627", x"0627", x"0628", x"0628", x"0628", x"0628", x"0629", x"0629", x"0629", x"0629", x"062a", x"062a", x"062a", x"062a", x"062b", x"062b", x"062b", x"062b", x"062c", x"062c", x"062c", x"062c", x"062c", x"062d", x"062d", x"062d", x"062d", x"062e", x"062e", x"062e", x"062e", x"062f", x"062f", x"062f", x"062f", x"0630", x"0630", x"0630", x"0630", x"0630", x"0631", x"0631", x"0631", x"0631", x"0632", x"0632", x"0632", x"0632", x"0633", x"0633", x"0633", x"0633", x"0634", x"0634", x"0634", x"0634", x"0635", x"0635", x"0635", x"0635", x"0635", x"0636", x"0636", x"0636", x"0636", x"0637", x"0637", x"0637", x"0637", x"0638", x"0638", x"0638", x"0638", x"0639", x"0639", x"0639", x"0639", x"063a", x"063a", x"063a", x"063a", x"063a", x"063b", x"063b", x"063b", x"063b", x"063c", x"063c", x"063c", x"063c", x"063d", x"063d", x"063d", x"063d", x"063e", x"063e", x"063e", x"063e", x"063e", x"063f", x"063f", x"063f", x"063f", x"0640", x"0640", x"0640", x"0640", x"0641", x"0641", x"0641", x"0641", x"0642", x"0642", x"0642", x"0642", x"0643", x"0643", x"0643", x"0643", x"0643", x"0644", x"0644", x"0644", x"0644", x"0645", x"0645", x"0645", x"0645", x"0646", x"0646", x"0646", x"0646", x"0647", x"0647", x"0647", x"0647", x"0648", x"0648", x"0648", x"0648", x"0649", x"0649", x"0649", x"0649", x"0649", x"064a", x"064a", x"064a", x"064a", x"064b", x"064b", x"064b", x"064b", x"064c", x"064c", x"064c", x"064c", x"064d", x"064d", x"064d", x"064d", x"064e", x"064e", x"064e", x"064e", x"064e", x"064f", x"064f", x"064f", x"064f", x"0650", x"0650", x"0650", x"0650", x"0651", x"0651", x"0651", x"0651", x"0652", x"0652", x"0652", x"0652", x"0653", x"0653", x"0653", x"0653", x"0653", x"0654", x"0654", x"0654", x"0654", x"0655", x"0655", x"0655", x"0655", x"0656", x"0656", x"0656", x"0656", x"0657", x"0657", x"0657", x"0657", x"0658", x"0658", x"0658", x"0658", x"0659", x"0659", x"0659", x"0659", x"0659", x"065a", x"065a", x"065a", x"065a", x"065b", x"065b", x"065b", x"065b", x"065c", x"065c", x"065c", x"065c", x"065d", x"065d", x"065d", x"065d", x"065e", x"065e", x"065e", x"065e", x"065e", x"065f", x"065f", x"065f", x"065f", x"0660", x"0660", x"0660", x"0660", x"0661", x"0661", x"0661", x"0661", x"0662", x"0662", x"0662", x"0662", x"0663", x"0663", x"0663", x"0663", x"0664", x"0664", x"0664", x"0664", x"0664", x"0665", x"0665", x"0665", x"0665", x"0666", x"0666", x"0666", x"0666", x"0667", x"0667", x"0667", x"0667", x"0668", x"0668", x"0668", x"0668", x"0669", x"0669", x"0669", x"0669", x"066a", x"066a", x"066a", x"066a", x"066a", x"066b", x"066b", x"066b", x"066b", x"066c", x"066c", x"066c", x"066c", x"066d", x"066d", x"066d", x"066d", x"066e", x"066e", x"066e", x"066e", x"066f", x"066f", x"066f", x"066f", x"0670", x"0670", x"0670", x"0670", x"0670", x"0671", x"0671", x"0671", x"0671", x"0672", x"0672", x"0672", x"0672", x"0673", x"0673", x"0673", x"0673", x"0674", x"0674", x"0674", x"0674", x"0675", x"0675", x"0675", x"0675", x"0676", x"0676", x"0676", x"0676", x"0677", x"0677", x"0677", x"0677", x"0677", x"0678", x"0678", x"0678", x"0678", x"0679", x"0679", x"0679", x"0679", x"067a", x"067a", x"067a", x"067a", x"067b", x"067b", x"067b", x"067b", x"067c", x"067c", x"067c", x"067c", x"067d", x"067d", x"067d", x"067d", x"067d", x"067e", x"067e", x"067e", x"067e", x"067f", x"067f", x"067f", x"067f", x"0680", x"0680", x"0680", x"0680", x"0681", x"0681", x"0681", x"0681", x"0682", x"0682", x"0682", x"0682", x"0683", x"0683", x"0683", x"0683", x"0684", x"0684", x"0684", x"0684", x"0684", x"0685", x"0685", x"0685", x"0685", x"0686", x"0686", x"0686", x"0686", x"0687", x"0687", x"0687", x"0687", x"0688", x"0688", x"0688", x"0688", x"0689", x"0689", x"0689", x"0689", x"068a", x"068a", x"068a", x"068a", x"068b", x"068b", x"068b", x"068b", x"068c", x"068c", x"068c", x"068c", x"068c", x"068d", x"068d", x"068d", x"068d", x"068e", x"068e", x"068e", x"068e", x"068f", x"068f", x"068f", x"068f", x"0690", x"0690", x"0690", x"0690", x"0691", x"0691", x"0691", x"0691", x"0692", x"0692", x"0692", x"0692", x"0693", x"0693", x"0693", x"0693", x"0693", x"0694", x"0694", x"0694", x"0694", x"0695", x"0695", x"0695", x"0695", x"0696", x"0696", x"0696", x"0696", x"0697", x"0697", x"0697", x"0697", x"0698", x"0698", x"0698", x"0698", x"0699", x"0699", x"0699", x"0699", x"069a", x"069a", x"069a", x"069a", x"069b", x"069b", x"069b", x"069b", x"069b", x"069c", x"069c", x"069c", x"069c", x"069d", x"069d", x"069d", x"069d", x"069e", x"069e", x"069e", x"069e", x"069f", x"069f", x"069f", x"069f", x"06a0", x"06a0", x"06a0", x"06a0", x"06a1", x"06a1", x"06a1", x"06a1", x"06a2", x"06a2", x"06a2", x"06a2", x"06a3", x"06a3", x"06a3", x"06a3", x"06a3", x"06a4", x"06a4", x"06a4", x"06a4", x"06a5", x"06a5", x"06a5", x"06a5", x"06a6", x"06a6", x"06a6", x"06a6", x"06a7", x"06a7", x"06a7", x"06a7", x"06a8", x"06a8", x"06a8", x"06a8", x"06a9", x"06a9", x"06a9", x"06a9", x"06aa", x"06aa", x"06aa", x"06aa", x"06ab", x"06ab", x"06ab", x"06ab", x"06ab", x"06ac", x"06ac", x"06ac", x"06ac", x"06ad", x"06ad", x"06ad", x"06ad", x"06ae", x"06ae", x"06ae", x"06ae", x"06af", x"06af", x"06af", x"06af", x"06b0", x"06b0", x"06b0", x"06b0", x"06b1", x"06b1", x"06b1", x"06b1", x"06b2", x"06b2", x"06b2", x"06b2", x"06b3", x"06b3", x"06b3", x"06b3", x"06b4", x"06b4", x"06b4", x"06b4", x"06b4", x"06b5", x"06b5", x"06b5", x"06b5", x"06b6", x"06b6", x"06b6", x"06b6", x"06b7", x"06b7", x"06b7", x"06b7", x"06b8", x"06b8", x"06b8", x"06b8", x"06b9", x"06b9", x"06b9", x"06b9", x"06ba", x"06ba", x"06ba", x"06ba", x"06bb", x"06bb", x"06bb", x"06bb", x"06bc", x"06bc", x"06bc", x"06bc", x"06bd", x"06bd", x"06bd", x"06bd", x"06be", x"06be", x"06be", x"06be", x"06be", x"06bf", x"06bf", x"06bf", x"06bf", x"06c0", x"06c0", x"06c0", x"06c0", x"06c1", x"06c1", x"06c1", x"06c1", x"06c2", x"06c2", x"06c2", x"06c2", x"06c3", x"06c3", x"06c3", x"06c3", x"06c4", x"06c4", x"06c4", x"06c4", x"06c5", x"06c5", x"06c5", x"06c5", x"06c6", x"06c6", x"06c6", x"06c6", x"06c7", x"06c7", x"06c7", x"06c7", x"06c8", x"06c8", x"06c8", x"06c8", x"06c8", x"06c9", x"06c9", x"06c9", x"06c9", x"06ca", x"06ca", x"06ca", x"06ca", x"06cb", x"06cb", x"06cb", x"06cb", x"06cc", x"06cc", x"06cc", x"06cc", x"06cd", x"06cd", x"06cd", x"06cd", x"06ce", x"06ce", x"06ce", x"06ce", x"06cf", x"06cf", x"06cf", x"06cf", x"06d0", x"06d0", x"06d0", x"06d0", x"06d1", x"06d1", x"06d1", x"06d1", x"06d2", x"06d2", x"06d2", x"06d2", x"06d3", x"06d3", x"06d3", x"06d3", x"06d3", x"06d4", x"06d4", x"06d4", x"06d4", x"06d5", x"06d5", x"06d5", x"06d5", x"06d6", x"06d6", x"06d6", x"06d6", x"06d7", x"06d7", x"06d7", x"06d7", x"06d8", x"06d8", x"06d8", x"06d8", x"06d9", x"06d9", x"06d9", x"06d9", x"06da", x"06da", x"06da", x"06da", x"06db", x"06db", x"06db", x"06db", x"06dc", x"06dc", x"06dc", x"06dc", x"06dd", x"06dd", x"06dd", x"06dd", x"06de", x"06de", x"06de", x"06de", x"06df", x"06df", x"06df", x"06df", x"06df", x"06e0", x"06e0", x"06e0", x"06e0", x"06e1", x"06e1", x"06e1", x"06e1", x"06e2", x"06e2", x"06e2", x"06e2", x"06e3", x"06e3", x"06e3", x"06e3", x"06e4", x"06e4", x"06e4", x"06e4", x"06e5", x"06e5", x"06e5", x"06e5", x"06e6", x"06e6", x"06e6", x"06e6", x"06e7", x"06e7", x"06e7", x"06e7", x"06e8", x"06e8", x"06e8", x"06e8", x"06e9", x"06e9", x"06e9", x"06e9", x"06ea", x"06ea", x"06ea", x"06ea", x"06eb", x"06eb", x"06eb", x"06eb", x"06eb", x"06ec", x"06ec", x"06ec", x"06ec", x"06ed", x"06ed", x"06ed", x"06ed", x"06ee", x"06ee", x"06ee", x"06ee", x"06ef", x"06ef", x"06ef", x"06ef", x"06f0", x"06f0", x"06f0", x"06f0", x"06f1", x"06f1", x"06f1", x"06f1", x"06f2", x"06f2", x"06f2", x"06f2", x"06f3", x"06f3", x"06f3", x"06f3", x"06f4", x"06f4", x"06f4", x"06f4", x"06f5", x"06f5", x"06f5", x"06f5", x"06f6", x"06f6", x"06f6", x"06f6", x"06f7", x"06f7", x"06f7", x"06f7", x"06f8", x"06f8", x"06f8", x"06f8", x"06f9", x"06f9", x"06f9", x"06f9", x"06fa", x"06fa", x"06fa", x"06fa", x"06fa", x"06fb", x"06fb", x"06fb", x"06fb", x"06fc", x"06fc", x"06fc", x"06fc", x"06fd", x"06fd", x"06fd", x"06fd", x"06fe", x"06fe", x"06fe", x"06fe", x"06ff", x"06ff", x"06ff", x"06ff", x"0700", x"0700", x"0700", x"0700", x"0701", x"0701", x"0701", x"0701", x"0702", x"0702", x"0702", x"0702", x"0703", x"0703", x"0703", x"0703", x"0704", x"0704", x"0704", x"0704", x"0705", x"0705", x"0705", x"0705", x"0706", x"0706", x"0706", x"0706", x"0707", x"0707", x"0707", x"0707", x"0708", x"0708", x"0708", x"0708", x"0709", x"0709", x"0709", x"0709", x"0709", x"070a", x"070a", x"070a", x"070a", x"070b", x"070b", x"070b", x"070b", x"070c", x"070c", x"070c", x"070c", x"070d", x"070d", x"070d", x"070d", x"070e", x"070e", x"070e", x"070e", x"070f", x"070f", x"070f", x"070f", x"0710", x"0710", x"0710", x"0710", x"0711", x"0711", x"0711", x"0711", x"0712", x"0712", x"0712", x"0712", x"0713", x"0713", x"0713", x"0713", x"0714", x"0714", x"0714", x"0714", x"0715", x"0715", x"0715", x"0715", x"0716", x"0716", x"0716", x"0716", x"0717", x"0717", x"0717", x"0717", x"0718", x"0718", x"0718", x"0718", x"0719", x"0719", x"0719", x"0719", x"071a", x"071a", x"071a", x"071a", x"071b", x"071b", x"071b", x"071b", x"071b", x"071c", x"071c", x"071c", x"071c", x"071d", x"071d", x"071d", x"071d", x"071e", x"071e", x"071e", x"071e", x"071f", x"071f", x"071f", x"071f", x"0720", x"0720", x"0720", x"0720", x"0721", x"0721", x"0721", x"0721", x"0722", x"0722", x"0722", x"0722", x"0723", x"0723", x"0723", x"0723", x"0724", x"0724", x"0724", x"0724", x"0725", x"0725", x"0725", x"0725", x"0726", x"0726", x"0726", x"0726", x"0727", x"0727", x"0727", x"0727", x"0728", x"0728", x"0728", x"0728", x"0729", x"0729", x"0729", x"0729", x"072a", x"072a", x"072a", x"072a", x"072b", x"072b", x"072b", x"072b", x"072c", x"072c", x"072c", x"072c", x"072d", x"072d", x"072d", x"072d", x"072e", x"072e", x"072e", x"072e", x"072f", x"072f", x"072f", x"072f", x"0730", x"0730", x"0730", x"0730", x"0731", x"0731", x"0731", x"0731", x"0731", x"0732", x"0732", x"0732", x"0732", x"0733", x"0733", x"0733", x"0733", x"0734", x"0734", x"0734", x"0734", x"0735", x"0735", x"0735", x"0735", x"0736", x"0736", x"0736", x"0736", x"0737", x"0737", x"0737", x"0737", x"0738", x"0738", x"0738", x"0738", x"0739", x"0739", x"0739", x"0739", x"073a", x"073a", x"073a", x"073a", x"073b", x"073b", x"073b", x"073b", x"073c", x"073c", x"073c", x"073c", x"073d", x"073d", x"073d", x"073d", x"073e", x"073e", x"073e", x"073e", x"073f", x"073f", x"073f", x"073f", x"0740", x"0740", x"0740", x"0740", x"0741", x"0741", x"0741", x"0741", x"0742", x"0742", x"0742", x"0742", x"0743", x"0743", x"0743", x"0743", x"0744", x"0744", x"0744", x"0744", x"0745", x"0745", x"0745", x"0745", x"0746", x"0746", x"0746", x"0746", x"0747", x"0747", x"0747", x"0747", x"0748", x"0748", x"0748", x"0748", x"0749", x"0749", x"0749", x"0749", x"074a", x"074a", x"074a", x"074a", x"074b", x"074b", x"074b", x"074b", x"074c", x"074c", x"074c", x"074c", x"074c", x"074d", x"074d", x"074d", x"074d", x"074e", x"074e", x"074e", x"074e", x"074f", x"074f", x"074f", x"074f", x"0750", x"0750", x"0750", x"0750", x"0751", x"0751", x"0751", x"0751", x"0752", x"0752", x"0752", x"0752", x"0753", x"0753", x"0753", x"0753", x"0754", x"0754", x"0754", x"0754", x"0755", x"0755", x"0755", x"0755", x"0756", x"0756", x"0756", x"0756", x"0757", x"0757", x"0757", x"0757", x"0758", x"0758", x"0758", x"0758", x"0759", x"0759", x"0759", x"0759", x"075a", x"075a", x"075a", x"075a", x"075b", x"075b", x"075b", x"075b", x"075c", x"075c", x"075c", x"075c", x"075d", x"075d", x"075d", x"075d", x"075e", x"075e", x"075e", x"075e", x"075f", x"075f", x"075f", x"075f", x"0760", x"0760", x"0760", x"0760", x"0761", x"0761", x"0761", x"0761", x"0762", x"0762", x"0762", x"0762", x"0763", x"0763", x"0763", x"0763", x"0764", x"0764", x"0764", x"0764", x"0765", x"0765", x"0765", x"0765", x"0766", x"0766", x"0766", x"0766", x"0767", x"0767", x"0767", x"0767", x"0768", x"0768", x"0768", x"0768", x"0769", x"0769", x"0769", x"0769", x"076a", x"076a", x"076a", x"076a", x"076b", x"076b", x"076b", x"076b", x"076c", x"076c", x"076c", x"076c", x"076d", x"076d", x"076d", x"076d", x"076e", x"076e", x"076e", x"076e", x"076f", x"076f", x"076f", x"076f", x"0770", x"0770", x"0770", x"0770", x"0771", x"0771", x"0771", x"0771", x"0772", x"0772", x"0772", x"0772", x"0773", x"0773", x"0773", x"0773", x"0774", x"0774", x"0774", x"0774", x"0774", x"0775", x"0775", x"0775", x"0775", x"0776", x"0776", x"0776", x"0776", x"0777", x"0777", x"0777", x"0777", x"0778", x"0778", x"0778", x"0778", x"0779", x"0779", x"0779", x"0779", x"077a", x"077a", x"077a", x"077a", x"077b", x"077b", x"077b", x"077b", x"077c", x"077c", x"077c", x"077c", x"077d", x"077d", x"077d", x"077d", x"077e", x"077e", x"077e", x"077e", x"077f", x"077f", x"077f", x"077f", x"0780", x"0780", x"0780", x"0780", x"0781", x"0781", x"0781", x"0781", x"0782", x"0782", x"0782", x"0782", x"0783", x"0783", x"0783", x"0783", x"0784", x"0784", x"0784", x"0784", x"0785", x"0785", x"0785", x"0785", x"0786", x"0786", x"0786", x"0786", x"0787", x"0787", x"0787", x"0787", x"0788", x"0788", x"0788", x"0788", x"0789", x"0789", x"0789", x"0789", x"078a", x"078a", x"078a", x"078a", x"078b", x"078b", x"078b", x"078b", x"078c", x"078c", x"078c", x"078c", x"078d", x"078d", x"078d", x"078d", x"078e", x"078e", x"078e", x"078e", x"078f", x"078f", x"078f", x"078f", x"0790", x"0790", x"0790", x"0790", x"0791", x"0791", x"0791", x"0791", x"0792", x"0792", x"0792", x"0792", x"0793", x"0793", x"0793", x"0793", x"0794", x"0794", x"0794", x"0794", x"0795", x"0795", x"0795", x"0795", x"0796", x"0796", x"0796", x"0796", x"0797", x"0797", x"0797", x"0797", x"0798", x"0798", x"0798", x"0798", x"0799", x"0799", x"0799", x"0799", x"079a", x"079a", x"079a", x"079a", x"079b", x"079b", x"079b", x"079b", x"079c", x"079c", x"079c", x"079c", x"079d", x"079d", x"079d", x"079d", x"079e", x"079e", x"079e", x"079e", x"079f", x"079f", x"079f", x"079f", x"07a0", x"07a0", x"07a0", x"07a0", x"07a1", x"07a1", x"07a1", x"07a1", x"07a2", x"07a2", x"07a2", x"07a2", x"07a3", x"07a3", x"07a3", x"07a3", x"07a4", x"07a4", x"07a4", x"07a4", x"07a5", x"07a5", x"07a5", x"07a5", x"07a6", x"07a6", x"07a6", x"07a6", x"07a7", x"07a7", x"07a7", x"07a7", x"07a8", x"07a8", x"07a8", x"07a8", x"07a9", x"07a9", x"07a9", x"07a9", x"07aa", x"07aa", x"07aa", x"07aa", x"07ab", x"07ab", x"07ab", x"07ab", x"07ac", x"07ac", x"07ac", x"07ac", x"07ad", x"07ad", x"07ad", x"07ad", x"07ae", x"07ae", x"07ae", x"07ae", x"07af", x"07af", x"07af", x"07af", x"07b0", x"07b0", x"07b0", x"07b0", x"07b1", x"07b1", x"07b1", x"07b1", x"07b2", x"07b2", x"07b2", x"07b2", x"07b3", x"07b3", x"07b3", x"07b3", x"07b4", x"07b4", x"07b4", x"07b4", x"07b5", x"07b5", x"07b5", x"07b5", x"07b6", x"07b6", x"07b6", x"07b6", x"07b7", x"07b7", x"07b7", x"07b7", x"07b8", x"07b8", x"07b8", x"07b8", x"07b9", x"07b9", x"07b9", x"07b9", x"07ba", x"07ba", x"07ba", x"07ba", x"07bb", x"07bb", x"07bb", x"07bb", x"07bc", x"07bc", x"07bc", x"07bc", x"07bd", x"07bd", x"07bd", x"07bd", x"07be", x"07be", x"07be", x"07be", x"07bf", x"07bf", x"07bf", x"07bf", x"07c0", x"07c0", x"07c0", x"07c0", x"07c1", x"07c1", x"07c1", x"07c1", x"07c2", x"07c2", x"07c2", x"07c2", x"07c3", x"07c3", x"07c3", x"07c3", x"07c4", x"07c4", x"07c4", x"07c4", x"07c5", x"07c5", x"07c5", x"07c5", x"07c6", x"07c6", x"07c6", x"07c6", x"07c7", x"07c7", x"07c7", x"07c7", x"07c8", x"07c8", x"07c8", x"07c8", x"07c9", x"07c9", x"07c9", x"07c9", x"07ca", x"07ca", x"07ca", x"07ca", x"07cb", x"07cb", x"07cb", x"07cb", x"07cc", x"07cc", x"07cc", x"07cc", x"07cd", x"07cd", x"07cd", x"07cd", x"07ce", x"07ce", x"07ce", x"07ce", x"07cf", x"07cf", x"07cf", x"07cf", x"07d0", x"07d0", x"07d0", x"07d0", x"07d1", x"07d1", x"07d1", x"07d1", x"07d2", x"07d2", x"07d2", x"07d2", x"07d3", x"07d3", x"07d3", x"07d3", x"07d4", x"07d4", x"07d4", x"07d4", x"07d5", x"07d5", x"07d5", x"07d5", x"07d6", x"07d6", x"07d6", x"07d6", x"07d7", x"07d7", x"07d7", x"07d7", x"07d8", x"07d8", x"07d8", x"07d8", x"07d9", x"07d9", x"07d9", x"07d9", x"07da", x"07da", x"07da", x"07da", x"07db", x"07db", x"07db", x"07db", x"07dc", x"07dc", x"07dc", x"07dc", x"07dd", x"07dd", x"07dd", x"07dd", x"07de", x"07de", x"07de", x"07de", x"07df", x"07df", x"07df", x"07df", x"07e0", x"07e0", x"07e0", x"07e0", x"07e1", x"07e1", x"07e1", x"07e1", x"07e2", x"07e2", x"07e2", x"07e2", x"07e3", x"07e3", x"07e3", x"07e3", x"07e4", x"07e4", x"07e4", x"07e4", x"07e5", x"07e5", x"07e5", x"07e5", x"07e6", x"07e6", x"07e6", x"07e6", x"07e7", x"07e7", x"07e7", x"07e7", x"07e8", x"07e8", x"07e8", x"07e8", x"07e9", x"07e9", x"07e9", x"07e9", x"07ea", x"07ea", x"07ea", x"07ea", x"07eb", x"07eb", x"07eb", x"07eb", x"07ec", x"07ec", x"07ec", x"07ec", x"07ed", x"07ed", x"07ed", x"07ed", x"07ee", x"07ee", x"07ee", x"07ee", x"07ef", x"07ef", x"07ef", x"07ef", x"07f0", x"07f0", x"07f0", x"07f0", x"07f1", x"07f1", x"07f1", x"07f1", x"07f2", x"07f2", x"07f2", x"07f2", x"07f3", x"07f3", x"07f3", x"07f3", x"07f4", x"07f4", x"07f4", x"07f4", x"07f5", x"07f5", x"07f5", x"07f5", x"07f6", x"07f6", x"07f6", x"07f6", x"07f7", x"07f7", x"07f7", x"07f7", x"07f8", x"07f8", x"07f8", x"07f8", x"07f9", x"07f9", x"07f9", x"07f9", x"07fa", x"07fa", x"07fa", x"07fa", x"07fb", x"07fb", x"07fb", x"07fb", x"07fc", x"07fc", x"07fc", x"07fc", x"07fd", x"07fd", x"07fd", x"07fd", x"07fe", x"07fe", x"07fe", x"07fe", x"07ff", x"07ff");
       begin

    process(Y)
    begin
	 O <= sigmoid_val(to_integer(unsigned(Y)));
    end process;

end Behavioral;

